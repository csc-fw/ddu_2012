//
// Design: incntrl
// Description: This top level Verilog model is created 
//              automatically by FusionHDL.
//

module Top;

defparam
 _7I5013_$1I4488_$1I4621.INIT_A = 9'H000,
 _7I5013_$1I4488_$1I4621.INIT_B = 18'H00000,
 _7I5013_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _7I5013_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _7I5013_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _7I5013_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _7I5013_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_A = 9'H000,
 _7I5013_$1I4488_$1I4620.INIT_B = 18'H00000,
 _7I5013_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _7I5013_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _7I5013_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _7I5013_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _7I5013_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I5013_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_A = 9'H000,
 _7I4974_$1I4488_$1I4621.INIT_B = 18'H00000,
 _7I4974_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _7I4974_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _7I4974_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _7I4974_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _7I4974_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_A = 9'H000,
 _7I4974_$1I4488_$1I4620.INIT_B = 18'H00000,
 _7I4974_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _7I4974_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _7I4974_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _7I4974_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _7I4974_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4974_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_A = 9'H000,
 _7I4863_$1I4488_$1I4621.INIT_B = 18'H00000,
 _7I4863_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _7I4863_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _7I4863_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _7I4863_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _7I4863_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_A = 9'H000,
 _7I4863_$1I4488_$1I4620.INIT_B = 18'H00000,
 _7I4863_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _7I4863_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _7I4863_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _7I4863_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _7I4863_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4863_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_A = 9'H000,
 _7I4838_$1I4488_$1I4621.INIT_B = 18'H00000,
 _7I4838_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _7I4838_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _7I4838_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _7I4838_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _7I4838_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_A = 9'H000,
 _7I4838_$1I4488_$1I4620.INIT_B = 18'H00000,
 _7I4838_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _7I4838_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _7I4838_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _7I4838_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _7I4838_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4838_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_A = 9'H000,
 _7I4762_$1I4488_$1I4621.INIT_B = 18'H00000,
 _7I4762_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _7I4762_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _7I4762_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _7I4762_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _7I4762_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_A = 9'H000,
 _7I4762_$1I4488_$1I4620.INIT_B = 18'H00000,
 _7I4762_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _7I4762_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _7I4762_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _7I4762_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _7I4762_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4762_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_A = 9'H000,
 _7I4731_$1I4488_$1I4621.INIT_B = 18'H00000,
 _7I4731_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _7I4731_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _7I4731_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _7I4731_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _7I4731_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_A = 9'H000,
 _7I4731_$1I4488_$1I4620.INIT_B = 18'H00000,
 _7I4731_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _7I4731_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _7I4731_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _7I4731_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _7I4731_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4731_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_A = 9'H000,
 _7I4712_$1I4488_$1I4621.INIT_B = 18'H00000,
 _7I4712_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _7I4712_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _7I4712_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _7I4712_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _7I4712_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_A = 9'H000,
 _7I4712_$1I4488_$1I4620.INIT_B = 18'H00000,
 _7I4712_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _7I4712_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _7I4712_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _7I4712_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _7I4712_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4712_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_A = 9'H000,
 _7I4651_$1I4488_$1I4621.INIT_B = 18'H00000,
 _7I4651_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _7I4651_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _7I4651_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _7I4651_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _7I4651_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_A = 9'H000,
 _7I4651_$1I4488_$1I4620.INIT_B = 18'H00000,
 _7I4651_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _7I4651_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _7I4651_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _7I4651_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _7I4651_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4651_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_A = 9'H000,
 _7I4632_$1I4488_$1I4621.INIT_B = 18'H00000,
 _7I4632_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _7I4632_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _7I4632_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _7I4632_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _7I4632_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_A = 9'H000,
 _7I4632_$1I4488_$1I4620.INIT_B = 18'H00000,
 _7I4632_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _7I4632_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _7I4632_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _7I4632_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _7I4632_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4632_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_A = 9'H000,
 _7I4616_$1I4488_$1I4621.INIT_B = 18'H00000,
 _7I4616_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _7I4616_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _7I4616_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _7I4616_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _7I4616_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_A = 9'H000,
 _7I4616_$1I4488_$1I4620.INIT_B = 18'H00000,
 _7I4616_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _7I4616_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _7I4616_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _7I4616_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _7I4616_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4616_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_A = 9'H000,
 _7I4615_$1I4488_$1I4621.INIT_B = 18'H00000,
 _7I4615_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _7I4615_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _7I4615_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _7I4615_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _7I4615_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_A = 9'H000,
 _7I4615_$1I4488_$1I4620.INIT_B = 18'H00000,
 _7I4615_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _7I4615_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _7I4615_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _7I4615_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _7I4615_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4615_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_A = 9'H000,
 _7I4614_$1I4488_$1I4621.INIT_B = 18'H00000,
 _7I4614_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _7I4614_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _7I4614_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _7I4614_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _7I4614_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_A = 9'H000,
 _7I4614_$1I4488_$1I4620.INIT_B = 18'H00000,
 _7I4614_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _7I4614_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _7I4614_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _7I4614_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _7I4614_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _7I4614_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_A = 9'H000,
 _6I4686_$1I4488_$1I4621.INIT_B = 18'H00000,
 _6I4686_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _6I4686_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _6I4686_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _6I4686_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _6I4686_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_A = 9'H000,
 _6I4686_$1I4488_$1I4620.INIT_B = 18'H00000,
 _6I4686_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _6I4686_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _6I4686_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _6I4686_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _6I4686_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4686_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_A = 9'H000,
 _6I4641_$1I4488_$1I4621.INIT_B = 18'H00000,
 _6I4641_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _6I4641_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _6I4641_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _6I4641_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _6I4641_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_A = 9'H000,
 _6I4641_$1I4488_$1I4620.INIT_B = 18'H00000,
 _6I4641_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _6I4641_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _6I4641_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _6I4641_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _6I4641_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4641_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_A = 9'H000,
 _6I4614_$1I4488_$1I4621.INIT_B = 18'H00000,
 _6I4614_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _6I4614_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _6I4614_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _6I4614_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _6I4614_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_A = 9'H000,
 _6I4614_$1I4488_$1I4620.INIT_B = 18'H00000,
 _6I4614_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _6I4614_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _6I4614_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _6I4614_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _6I4614_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4614_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_A = 9'H000,
 _6I4598_$1I4488_$1I4621.INIT_B = 18'H00000,
 _6I4598_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _6I4598_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _6I4598_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _6I4598_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _6I4598_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_A = 9'H000,
 _6I4598_$1I4488_$1I4620.INIT_B = 18'H00000,
 _6I4598_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _6I4598_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _6I4598_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _6I4598_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _6I4598_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4598_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_A = 9'H000,
 _6I4575_$1I4488_$1I4621.INIT_B = 18'H00000,
 _6I4575_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _6I4575_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _6I4575_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _6I4575_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _6I4575_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_A = 9'H000,
 _6I4575_$1I4488_$1I4620.INIT_B = 18'H00000,
 _6I4575_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _6I4575_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _6I4575_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _6I4575_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _6I4575_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4575_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_A = 9'H000,
 _6I4529_$1I4488_$1I4621.INIT_B = 18'H00000,
 _6I4529_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _6I4529_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _6I4529_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _6I4529_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _6I4529_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_A = 9'H000,
 _6I4529_$1I4488_$1I4620.INIT_B = 18'H00000,
 _6I4529_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _6I4529_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _6I4529_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _6I4529_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _6I4529_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4529_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_A = 9'H000,
 _6I4504_$1I4488_$1I4621.INIT_B = 18'H00000,
 _6I4504_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _6I4504_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _6I4504_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _6I4504_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _6I4504_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_A = 9'H000,
 _6I4504_$1I4488_$1I4620.INIT_B = 18'H00000,
 _6I4504_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _6I4504_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _6I4504_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _6I4504_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _6I4504_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4504_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_A = 9'H000,
 _6I4479_$1I4488_$1I4621.INIT_B = 18'H00000,
 _6I4479_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _6I4479_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _6I4479_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _6I4479_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _6I4479_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_A = 9'H000,
 _6I4479_$1I4488_$1I4620.INIT_B = 18'H00000,
 _6I4479_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _6I4479_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _6I4479_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _6I4479_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _6I4479_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4479_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4446_$1I3863.ALIGN_COMMA_MSB = TRUE,
 _6I4446_$1I3863.CHAN_BOND_LIMIT = 16,
 _6I4446_$1I3863.CHAN_BOND_MODE = "OFF",
 _6I4446_$1I3863.CHAN_BOND_OFFSET = 8,
 _6I4446_$1I3863.CHAN_BOND_ONE_SHOT = "FALSE",
 _6I4446_$1I3863.CHAN_BOND_SEQ_1_1 = 11'B00000000000,
 _6I4446_$1I3863.CHAN_BOND_SEQ_1_2 = 11'B00000000000,
 _6I4446_$1I3863.CHAN_BOND_SEQ_1_3 = 11'B00000000000,
 _6I4446_$1I3863.CHAN_BOND_SEQ_1_4 = 11'B00000000000,
 _6I4446_$1I3863.CHAN_BOND_SEQ_2_1 = 11'B00000000000,
 _6I4446_$1I3863.CHAN_BOND_SEQ_2_2 = 11'B00000000000,
 _6I4446_$1I3863.CHAN_BOND_SEQ_2_3 = 11'B00000000000,
 _6I4446_$1I3863.CHAN_BOND_SEQ_2_4 = 11'B00000000000,
 _6I4446_$1I3863.CHAN_BOND_SEQ_2_USE = "FALSE",
 _6I4446_$1I3863.CHAN_BOND_SEQ_LEN = 1,
 _6I4446_$1I3863.CHAN_BOND_WAIT = 8,
 _6I4446_$1I3863.CLK_COR_INSERT_IDLE_FLAG = "FALSE",
 _6I4446_$1I3863.CLK_COR_KEEP_IDLE = TRUE,
 _6I4446_$1I3863.CLK_COR_REPEAT_WAIT = 0,
 _6I4446_$1I3863.CLK_COR_SEQ_1_1 = 00110111100,
 _6I4446_$1I3863.CLK_COR_SEQ_1_2 = 00011000101,
 _6I4446_$1I3863.CLK_COR_SEQ_1_3 = 11'B00000000000,
 _6I4446_$1I3863.CLK_COR_SEQ_1_4 = 11'B00000000000,
 _6I4446_$1I3863.CLK_COR_SEQ_2_1 = 00110111100,
 _6I4446_$1I3863.CLK_COR_SEQ_2_2 = 00001010000,
 _6I4446_$1I3863.CLK_COR_SEQ_2_3 = 11'B00000000000,
 _6I4446_$1I3863.CLK_COR_SEQ_2_4 = 11'B00000000000,
 _6I4446_$1I3863.CLK_COR_SEQ_2_USE = TRUE,
 _6I4446_$1I3863.CLK_COR_SEQ_LEN = 2,
 _6I4446_$1I3863.CLK_CORRECT_USE = "TRUE",
 _6I4446_$1I3863.COMMA_10B_MASK = 10'B1111111000,
 _6I4446_$1I3863.CRC_END_OF_PKT = "K29_7",
 _6I4446_$1I3863.CRC_FORMAT = "USER_MODE",
 _6I4446_$1I3863.CRC_START_OF_PKT = "K27_7",
 _6I4446_$1I3863.DEC_MCOMMA_DETECT = "TRUE",
 _6I4446_$1I3863.DEC_PCOMMA_DETECT = "TRUE",
 _6I4446_$1I3863.DEC_VALID_COMMA_ONLY = "TRUE",
 _6I4446_$1I3863.MCOMMA_10B_VALUE = 10'B1100000000,
 _6I4446_$1I3863.MCOMMA_DETECT = "TRUE",
 _6I4446_$1I3863.PCOMMA_10B_VALUE = 10'B0011111000,
 _6I4446_$1I3863.PCOMMA_DETECT = "TRUE",
 _6I4446_$1I3863.REF_CLK_V_SEL = 1,
 _6I4446_$1I3863.RX_BUFFER_USE = "TRUE",
 _6I4446_$1I3863.RX_CRC_USE = "FALSE",
 _6I4446_$1I3863.RX_DATA_WIDTH = 2,
 _6I4446_$1I3863.RX_DECODE_USE = "TRUE",
 _6I4446_$1I3863.RX_LOS_INVALID_INCR = 2,
 _6I4446_$1I3863.RX_LOS_THRESHOLD = 8,
 _6I4446_$1I3863.RX_LOSS_OF_SYNC_FSM = "TRUE",
 _6I4446_$1I3863.SERDES_10B = "FALSE",
 _6I4446_$1I3863.TERMINATION_IMP = 50,
 _6I4446_$1I3863.TX_BUFFER_USE = "TRUE",
 _6I4446_$1I3863.TX_CRC_FORCE_VALUE = 8'B11010110,
 _6I4446_$1I3863.TX_CRC_USE = "FALSE",
 _6I4446_$1I3863.TX_DATA_WIDTH = 2,
 _6I4446_$1I3863.TX_DIFF_CTRL = 400,
 _6I4446_$1I3863.TX_PREEMPHASIS = 0,
 _6I4415_$1I3863.ALIGN_COMMA_MSB = TRUE,
 _6I4415_$1I3863.CHAN_BOND_LIMIT = 16,
 _6I4415_$1I3863.CHAN_BOND_MODE = "OFF",
 _6I4415_$1I3863.CHAN_BOND_OFFSET = 8,
 _6I4415_$1I3863.CHAN_BOND_ONE_SHOT = "FALSE",
 _6I4415_$1I3863.CHAN_BOND_SEQ_1_1 = 11'B00000000000,
 _6I4415_$1I3863.CHAN_BOND_SEQ_1_2 = 11'B00000000000,
 _6I4415_$1I3863.CHAN_BOND_SEQ_1_3 = 11'B00000000000,
 _6I4415_$1I3863.CHAN_BOND_SEQ_1_4 = 11'B00000000000,
 _6I4415_$1I3863.CHAN_BOND_SEQ_2_1 = 11'B00000000000,
 _6I4415_$1I3863.CHAN_BOND_SEQ_2_2 = 11'B00000000000,
 _6I4415_$1I3863.CHAN_BOND_SEQ_2_3 = 11'B00000000000,
 _6I4415_$1I3863.CHAN_BOND_SEQ_2_4 = 11'B00000000000,
 _6I4415_$1I3863.CHAN_BOND_SEQ_2_USE = "FALSE",
 _6I4415_$1I3863.CHAN_BOND_SEQ_LEN = 1,
 _6I4415_$1I3863.CHAN_BOND_WAIT = 8,
 _6I4415_$1I3863.CLK_COR_INSERT_IDLE_FLAG = "FALSE",
 _6I4415_$1I3863.CLK_COR_KEEP_IDLE = TRUE,
 _6I4415_$1I3863.CLK_COR_REPEAT_WAIT = 0,
 _6I4415_$1I3863.CLK_COR_SEQ_1_1 = 00110111100,
 _6I4415_$1I3863.CLK_COR_SEQ_1_2 = 00011000101,
 _6I4415_$1I3863.CLK_COR_SEQ_1_3 = 11'B00000000000,
 _6I4415_$1I3863.CLK_COR_SEQ_1_4 = 11'B00000000000,
 _6I4415_$1I3863.CLK_COR_SEQ_2_1 = 00110111100,
 _6I4415_$1I3863.CLK_COR_SEQ_2_2 = 00001010000,
 _6I4415_$1I3863.CLK_COR_SEQ_2_3 = 11'B00000000000,
 _6I4415_$1I3863.CLK_COR_SEQ_2_4 = 11'B00000000000,
 _6I4415_$1I3863.CLK_COR_SEQ_2_USE = TRUE,
 _6I4415_$1I3863.CLK_COR_SEQ_LEN = 2,
 _6I4415_$1I3863.CLK_CORRECT_USE = "TRUE",
 _6I4415_$1I3863.COMMA_10B_MASK = 10'B1111111000,
 _6I4415_$1I3863.CRC_END_OF_PKT = "K29_7",
 _6I4415_$1I3863.CRC_FORMAT = "USER_MODE",
 _6I4415_$1I3863.CRC_START_OF_PKT = "K27_7",
 _6I4415_$1I3863.DEC_MCOMMA_DETECT = "TRUE",
 _6I4415_$1I3863.DEC_PCOMMA_DETECT = "TRUE",
 _6I4415_$1I3863.DEC_VALID_COMMA_ONLY = "TRUE",
 _6I4415_$1I3863.MCOMMA_10B_VALUE = 10'B1100000000,
 _6I4415_$1I3863.MCOMMA_DETECT = "TRUE",
 _6I4415_$1I3863.PCOMMA_10B_VALUE = 10'B0011111000,
 _6I4415_$1I3863.PCOMMA_DETECT = "TRUE",
 _6I4415_$1I3863.REF_CLK_V_SEL = 1,
 _6I4415_$1I3863.RX_BUFFER_USE = "TRUE",
 _6I4415_$1I3863.RX_CRC_USE = "FALSE",
 _6I4415_$1I3863.RX_DATA_WIDTH = 2,
 _6I4415_$1I3863.RX_DECODE_USE = "TRUE",
 _6I4415_$1I3863.RX_LOS_INVALID_INCR = 2,
 _6I4415_$1I3863.RX_LOS_THRESHOLD = 8,
 _6I4415_$1I3863.RX_LOSS_OF_SYNC_FSM = "TRUE",
 _6I4415_$1I3863.SERDES_10B = "FALSE",
 _6I4415_$1I3863.TERMINATION_IMP = 50,
 _6I4415_$1I3863.TX_BUFFER_USE = "TRUE",
 _6I4415_$1I3863.TX_CRC_FORCE_VALUE = 8'B11010110,
 _6I4415_$1I3863.TX_CRC_USE = "FALSE",
 _6I4415_$1I3863.TX_DATA_WIDTH = 2,
 _6I4415_$1I3863.TX_DIFF_CTRL = 400,
 _6I4415_$1I3863.TX_PREEMPHASIS = 0,
 _6I4412_$1I3863.ALIGN_COMMA_MSB = TRUE,
 _6I4412_$1I3863.CHAN_BOND_LIMIT = 16,
 _6I4412_$1I3863.CHAN_BOND_MODE = "OFF",
 _6I4412_$1I3863.CHAN_BOND_OFFSET = 8,
 _6I4412_$1I3863.CHAN_BOND_ONE_SHOT = "FALSE",
 _6I4412_$1I3863.CHAN_BOND_SEQ_1_1 = 11'B00000000000,
 _6I4412_$1I3863.CHAN_BOND_SEQ_1_2 = 11'B00000000000,
 _6I4412_$1I3863.CHAN_BOND_SEQ_1_3 = 11'B00000000000,
 _6I4412_$1I3863.CHAN_BOND_SEQ_1_4 = 11'B00000000000,
 _6I4412_$1I3863.CHAN_BOND_SEQ_2_1 = 11'B00000000000,
 _6I4412_$1I3863.CHAN_BOND_SEQ_2_2 = 11'B00000000000,
 _6I4412_$1I3863.CHAN_BOND_SEQ_2_3 = 11'B00000000000,
 _6I4412_$1I3863.CHAN_BOND_SEQ_2_4 = 11'B00000000000,
 _6I4412_$1I3863.CHAN_BOND_SEQ_2_USE = "FALSE",
 _6I4412_$1I3863.CHAN_BOND_SEQ_LEN = 1,
 _6I4412_$1I3863.CHAN_BOND_WAIT = 8,
 _6I4412_$1I3863.CLK_COR_INSERT_IDLE_FLAG = "FALSE",
 _6I4412_$1I3863.CLK_COR_KEEP_IDLE = TRUE,
 _6I4412_$1I3863.CLK_COR_REPEAT_WAIT = 0,
 _6I4412_$1I3863.CLK_COR_SEQ_1_1 = 00110111100,
 _6I4412_$1I3863.CLK_COR_SEQ_1_2 = 00011000101,
 _6I4412_$1I3863.CLK_COR_SEQ_1_3 = 11'B00000000000,
 _6I4412_$1I3863.CLK_COR_SEQ_1_4 = 11'B00000000000,
 _6I4412_$1I3863.CLK_COR_SEQ_2_1 = 00110111100,
 _6I4412_$1I3863.CLK_COR_SEQ_2_2 = 00001010000,
 _6I4412_$1I3863.CLK_COR_SEQ_2_3 = 11'B00000000000,
 _6I4412_$1I3863.CLK_COR_SEQ_2_4 = 11'B00000000000,
 _6I4412_$1I3863.CLK_COR_SEQ_2_USE = TRUE,
 _6I4412_$1I3863.CLK_COR_SEQ_LEN = 2,
 _6I4412_$1I3863.CLK_CORRECT_USE = "TRUE",
 _6I4412_$1I3863.COMMA_10B_MASK = 10'B1111111000,
 _6I4412_$1I3863.CRC_END_OF_PKT = "K29_7",
 _6I4412_$1I3863.CRC_FORMAT = "USER_MODE",
 _6I4412_$1I3863.CRC_START_OF_PKT = "K27_7",
 _6I4412_$1I3863.DEC_MCOMMA_DETECT = "TRUE",
 _6I4412_$1I3863.DEC_PCOMMA_DETECT = "TRUE",
 _6I4412_$1I3863.DEC_VALID_COMMA_ONLY = "TRUE",
 _6I4412_$1I3863.MCOMMA_10B_VALUE = 10'B1100000000,
 _6I4412_$1I3863.MCOMMA_DETECT = "TRUE",
 _6I4412_$1I3863.PCOMMA_10B_VALUE = 10'B0011111000,
 _6I4412_$1I3863.PCOMMA_DETECT = "TRUE",
 _6I4412_$1I3863.REF_CLK_V_SEL = 1,
 _6I4412_$1I3863.RX_BUFFER_USE = "TRUE",
 _6I4412_$1I3863.RX_CRC_USE = "FALSE",
 _6I4412_$1I3863.RX_DATA_WIDTH = 2,
 _6I4412_$1I3863.RX_DECODE_USE = "TRUE",
 _6I4412_$1I3863.RX_LOS_INVALID_INCR = 2,
 _6I4412_$1I3863.RX_LOS_THRESHOLD = 8,
 _6I4412_$1I3863.RX_LOSS_OF_SYNC_FSM = "TRUE",
 _6I4412_$1I3863.SERDES_10B = "FALSE",
 _6I4412_$1I3863.TERMINATION_IMP = 50,
 _6I4412_$1I3863.TX_BUFFER_USE = "TRUE",
 _6I4412_$1I3863.TX_CRC_FORCE_VALUE = 8'B11010110,
 _6I4412_$1I3863.TX_CRC_USE = "FALSE",
 _6I4412_$1I3863.TX_DATA_WIDTH = 2,
 _6I4412_$1I3863.TX_DIFF_CTRL = 400,
 _6I4412_$1I3863.TX_PREEMPHASIS = 0,
 _6I4143_$1I4488_$1I4621.INIT_A = 9'H000,
 _6I4143_$1I4488_$1I4621.INIT_B = 18'H00000,
 _6I4143_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _6I4143_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _6I4143_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _6I4143_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _6I4143_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_A = 9'H000,
 _6I4143_$1I4488_$1I4620.INIT_B = 18'H00000,
 _6I4143_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _6I4143_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _6I4143_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _6I4143_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _6I4143_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _6I4143_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4382_$1I3863.ALIGN_COMMA_MSB = TRUE,
 _5I4382_$1I3863.CHAN_BOND_LIMIT = 16,
 _5I4382_$1I3863.CHAN_BOND_MODE = "OFF",
 _5I4382_$1I3863.CHAN_BOND_OFFSET = 8,
 _5I4382_$1I3863.CHAN_BOND_ONE_SHOT = "FALSE",
 _5I4382_$1I3863.CHAN_BOND_SEQ_1_1 = 11'B00000000000,
 _5I4382_$1I3863.CHAN_BOND_SEQ_1_2 = 11'B00000000000,
 _5I4382_$1I3863.CHAN_BOND_SEQ_1_3 = 11'B00000000000,
 _5I4382_$1I3863.CHAN_BOND_SEQ_1_4 = 11'B00000000000,
 _5I4382_$1I3863.CHAN_BOND_SEQ_2_1 = 11'B00000000000,
 _5I4382_$1I3863.CHAN_BOND_SEQ_2_2 = 11'B00000000000,
 _5I4382_$1I3863.CHAN_BOND_SEQ_2_3 = 11'B00000000000,
 _5I4382_$1I3863.CHAN_BOND_SEQ_2_4 = 11'B00000000000,
 _5I4382_$1I3863.CHAN_BOND_SEQ_2_USE = "FALSE",
 _5I4382_$1I3863.CHAN_BOND_SEQ_LEN = 1,
 _5I4382_$1I3863.CHAN_BOND_WAIT = 8,
 _5I4382_$1I3863.CLK_COR_INSERT_IDLE_FLAG = "FALSE",
 _5I4382_$1I3863.CLK_COR_KEEP_IDLE = TRUE,
 _5I4382_$1I3863.CLK_COR_REPEAT_WAIT = 0,
 _5I4382_$1I3863.CLK_COR_SEQ_1_1 = 00110111100,
 _5I4382_$1I3863.CLK_COR_SEQ_1_2 = 00011000101,
 _5I4382_$1I3863.CLK_COR_SEQ_1_3 = 11'B00000000000,
 _5I4382_$1I3863.CLK_COR_SEQ_1_4 = 11'B00000000000,
 _5I4382_$1I3863.CLK_COR_SEQ_2_1 = 00110111100,
 _5I4382_$1I3863.CLK_COR_SEQ_2_2 = 00001010000,
 _5I4382_$1I3863.CLK_COR_SEQ_2_3 = 11'B00000000000,
 _5I4382_$1I3863.CLK_COR_SEQ_2_4 = 11'B00000000000,
 _5I4382_$1I3863.CLK_COR_SEQ_2_USE = TRUE,
 _5I4382_$1I3863.CLK_COR_SEQ_LEN = 2,
 _5I4382_$1I3863.CLK_CORRECT_USE = "TRUE",
 _5I4382_$1I3863.COMMA_10B_MASK = 10'B1111111000,
 _5I4382_$1I3863.CRC_END_OF_PKT = "K29_7",
 _5I4382_$1I3863.CRC_FORMAT = "USER_MODE",
 _5I4382_$1I3863.CRC_START_OF_PKT = "K27_7",
 _5I4382_$1I3863.DEC_MCOMMA_DETECT = "TRUE",
 _5I4382_$1I3863.DEC_PCOMMA_DETECT = "TRUE",
 _5I4382_$1I3863.DEC_VALID_COMMA_ONLY = "TRUE",
 _5I4382_$1I3863.MCOMMA_10B_VALUE = 10'B1100000000,
 _5I4382_$1I3863.MCOMMA_DETECT = "TRUE",
 _5I4382_$1I3863.PCOMMA_10B_VALUE = 10'B0011111000,
 _5I4382_$1I3863.PCOMMA_DETECT = "TRUE",
 _5I4382_$1I3863.REF_CLK_V_SEL = 1,
 _5I4382_$1I3863.RX_BUFFER_USE = "TRUE",
 _5I4382_$1I3863.RX_CRC_USE = "FALSE",
 _5I4382_$1I3863.RX_DATA_WIDTH = 2,
 _5I4382_$1I3863.RX_DECODE_USE = "TRUE",
 _5I4382_$1I3863.RX_LOS_INVALID_INCR = 2,
 _5I4382_$1I3863.RX_LOS_THRESHOLD = 8,
 _5I4382_$1I3863.RX_LOSS_OF_SYNC_FSM = "TRUE",
 _5I4382_$1I3863.SERDES_10B = "FALSE",
 _5I4382_$1I3863.TERMINATION_IMP = 50,
 _5I4382_$1I3863.TX_BUFFER_USE = "TRUE",
 _5I4382_$1I3863.TX_CRC_FORCE_VALUE = 8'B11010110,
 _5I4382_$1I3863.TX_CRC_USE = "FALSE",
 _5I4382_$1I3863.TX_DATA_WIDTH = 2,
 _5I4382_$1I3863.TX_DIFF_CTRL = 400,
 _5I4382_$1I3863.TX_PREEMPHASIS = 0,
 _5I4143_$1I4488_$1I4621.INIT_A = 9'H000,
 _5I4143_$1I4488_$1I4621.INIT_B = 18'H00000,
 _5I4143_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _5I4143_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _5I4143_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _5I4143_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _5I4143_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_A = 9'H000,
 _5I4143_$1I4488_$1I4620.INIT_B = 18'H00000,
 _5I4143_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _5I4143_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _5I4143_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _5I4143_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _5I4143_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _5I4143_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_A = 9'H000,
 _4I4657_$1I4488_$1I4621.INIT_B = 18'H00000,
 _4I4657_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _4I4657_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _4I4657_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _4I4657_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _4I4657_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_A = 9'H000,
 _4I4657_$1I4488_$1I4620.INIT_B = 18'H00000,
 _4I4657_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _4I4657_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _4I4657_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _4I4657_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _4I4657_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4657_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_A = 9'H000,
 _4I4630_$1I4488_$1I4621.INIT_B = 18'H00000,
 _4I4630_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _4I4630_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _4I4630_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _4I4630_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _4I4630_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_A = 9'H000,
 _4I4630_$1I4488_$1I4620.INIT_B = 18'H00000,
 _4I4630_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _4I4630_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _4I4630_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _4I4630_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _4I4630_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4630_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_A = 9'H000,
 _4I4611_$1I4488_$1I4621.INIT_B = 18'H00000,
 _4I4611_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _4I4611_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _4I4611_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _4I4611_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _4I4611_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_A = 9'H000,
 _4I4611_$1I4488_$1I4620.INIT_B = 18'H00000,
 _4I4611_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _4I4611_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _4I4611_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _4I4611_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _4I4611_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4611_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_A = 9'H000,
 _4I4560_$1I4488_$1I4621.INIT_B = 18'H00000,
 _4I4560_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _4I4560_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _4I4560_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _4I4560_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _4I4560_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_A = 9'H000,
 _4I4560_$1I4488_$1I4620.INIT_B = 18'H00000,
 _4I4560_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _4I4560_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _4I4560_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _4I4560_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _4I4560_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4560_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_A = 9'H000,
 _4I4526_$1I4488_$1I4621.INIT_B = 18'H00000,
 _4I4526_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _4I4526_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _4I4526_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _4I4526_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _4I4526_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_A = 9'H000,
 _4I4526_$1I4488_$1I4620.INIT_B = 18'H00000,
 _4I4526_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _4I4526_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _4I4526_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _4I4526_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _4I4526_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4526_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_A = 9'H000,
 _4I4501_$1I4488_$1I4621.INIT_B = 18'H00000,
 _4I4501_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _4I4501_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _4I4501_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _4I4501_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _4I4501_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_A = 9'H000,
 _4I4501_$1I4488_$1I4620.INIT_B = 18'H00000,
 _4I4501_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _4I4501_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _4I4501_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _4I4501_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _4I4501_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4501_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_A = 9'H000,
 _4I4476_$1I4488_$1I4621.INIT_B = 18'H00000,
 _4I4476_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _4I4476_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _4I4476_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _4I4476_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _4I4476_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_A = 9'H000,
 _4I4476_$1I4488_$1I4620.INIT_B = 18'H00000,
 _4I4476_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _4I4476_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _4I4476_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _4I4476_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _4I4476_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4476_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_A = 9'H000,
 _4I4475_$1I4488_$1I4621.INIT_B = 18'H00000,
 _4I4475_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _4I4475_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _4I4475_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _4I4475_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _4I4475_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_A = 9'H000,
 _4I4475_$1I4488_$1I4620.INIT_B = 18'H00000,
 _4I4475_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _4I4475_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _4I4475_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _4I4475_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _4I4475_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4475_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_A = 9'H000,
 _4I4426_$1I4488_$1I4621.INIT_B = 18'H00000,
 _4I4426_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _4I4426_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _4I4426_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _4I4426_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _4I4426_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_A = 9'H000,
 _4I4426_$1I4488_$1I4620.INIT_B = 18'H00000,
 _4I4426_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _4I4426_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _4I4426_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _4I4426_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _4I4426_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4426_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_A = 9'H000,
 _4I4399_$1I4488_$1I4621.INIT_B = 18'H00000,
 _4I4399_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _4I4399_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _4I4399_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _4I4399_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _4I4399_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_A = 9'H000,
 _4I4399_$1I4488_$1I4620.INIT_B = 18'H00000,
 _4I4399_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _4I4399_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _4I4399_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _4I4399_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _4I4399_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4399_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_A = 9'H000,
 _4I4365_$1I4488_$1I4621.INIT_B = 18'H00000,
 _4I4365_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _4I4365_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _4I4365_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _4I4365_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _4I4365_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_A = 9'H000,
 _4I4365_$1I4488_$1I4620.INIT_B = 18'H00000,
 _4I4365_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _4I4365_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _4I4365_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _4I4365_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _4I4365_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4365_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_A = 9'H000,
 _4I4329_$1I4488_$1I4621.INIT_B = 18'H00000,
 _4I4329_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _4I4329_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _4I4329_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _4I4329_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _4I4329_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_A = 9'H000,
 _4I4329_$1I4488_$1I4620.INIT_B = 18'H00000,
 _4I4329_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _4I4329_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _4I4329_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _4I4329_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _4I4329_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _4I4329_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_A = 9'H000,
 _3I4551_$1I4488_$1I4621.INIT_B = 18'H00000,
 _3I4551_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _3I4551_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _3I4551_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _3I4551_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _3I4551_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_A = 9'H000,
 _3I4551_$1I4488_$1I4620.INIT_B = 18'H00000,
 _3I4551_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _3I4551_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _3I4551_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _3I4551_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _3I4551_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4551_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_A = 9'H000,
 _3I4526_$1I4488_$1I4621.INIT_B = 18'H00000,
 _3I4526_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _3I4526_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _3I4526_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _3I4526_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _3I4526_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_A = 9'H000,
 _3I4526_$1I4488_$1I4620.INIT_B = 18'H00000,
 _3I4526_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _3I4526_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _3I4526_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _3I4526_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _3I4526_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4526_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_A = 9'H000,
 _3I4496_$1I4488_$1I4621.INIT_B = 18'H00000,
 _3I4496_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _3I4496_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _3I4496_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _3I4496_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _3I4496_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_A = 9'H000,
 _3I4496_$1I4488_$1I4620.INIT_B = 18'H00000,
 _3I4496_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _3I4496_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _3I4496_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _3I4496_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _3I4496_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4496_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_A = 9'H000,
 _3I4489_$1I4488_$1I4621.INIT_B = 18'H00000,
 _3I4489_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _3I4489_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _3I4489_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _3I4489_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _3I4489_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_A = 9'H000,
 _3I4489_$1I4488_$1I4620.INIT_B = 18'H00000,
 _3I4489_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _3I4489_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _3I4489_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _3I4489_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _3I4489_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4489_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_A = 9'H000,
 _3I4464_$1I4488_$1I4621.INIT_B = 18'H00000,
 _3I4464_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _3I4464_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _3I4464_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _3I4464_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _3I4464_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_A = 9'H000,
 _3I4464_$1I4488_$1I4620.INIT_B = 18'H00000,
 _3I4464_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _3I4464_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _3I4464_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _3I4464_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _3I4464_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4464_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_A = 9'H000,
 _3I4417_$1I4488_$1I4621.INIT_B = 18'H00000,
 _3I4417_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _3I4417_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _3I4417_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _3I4417_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _3I4417_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_A = 9'H000,
 _3I4417_$1I4488_$1I4620.INIT_B = 18'H00000,
 _3I4417_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _3I4417_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _3I4417_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _3I4417_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _3I4417_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4417_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_A = 9'H000,
 _3I4392_$1I4488_$1I4621.INIT_B = 18'H00000,
 _3I4392_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _3I4392_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _3I4392_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _3I4392_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _3I4392_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_A = 9'H000,
 _3I4392_$1I4488_$1I4620.INIT_B = 18'H00000,
 _3I4392_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _3I4392_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _3I4392_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _3I4392_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _3I4392_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4392_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_A = 9'H000,
 _3I4365_$1I4488_$1I4621.INIT_B = 18'H00000,
 _3I4365_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _3I4365_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _3I4365_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _3I4365_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _3I4365_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_A = 9'H000,
 _3I4365_$1I4488_$1I4620.INIT_B = 18'H00000,
 _3I4365_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _3I4365_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _3I4365_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _3I4365_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _3I4365_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4365_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_A = 9'H000,
 _3I4329_$1I4488_$1I4621.INIT_B = 18'H00000,
 _3I4329_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _3I4329_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _3I4329_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _3I4329_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _3I4329_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_A = 9'H000,
 _3I4329_$1I4488_$1I4620.INIT_B = 18'H00000,
 _3I4329_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _3I4329_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _3I4329_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _3I4329_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _3I4329_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4329_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _3I4274_$1I3863.ALIGN_COMMA_MSB = TRUE,
 _3I4274_$1I3863.CHAN_BOND_LIMIT = 16,
 _3I4274_$1I3863.CHAN_BOND_MODE = "OFF",
 _3I4274_$1I3863.CHAN_BOND_OFFSET = 8,
 _3I4274_$1I3863.CHAN_BOND_ONE_SHOT = "FALSE",
 _3I4274_$1I3863.CHAN_BOND_SEQ_1_1 = 11'B00000000000,
 _3I4274_$1I3863.CHAN_BOND_SEQ_1_2 = 11'B00000000000,
 _3I4274_$1I3863.CHAN_BOND_SEQ_1_3 = 11'B00000000000,
 _3I4274_$1I3863.CHAN_BOND_SEQ_1_4 = 11'B00000000000,
 _3I4274_$1I3863.CHAN_BOND_SEQ_2_1 = 11'B00000000000,
 _3I4274_$1I3863.CHAN_BOND_SEQ_2_2 = 11'B00000000000,
 _3I4274_$1I3863.CHAN_BOND_SEQ_2_3 = 11'B00000000000,
 _3I4274_$1I3863.CHAN_BOND_SEQ_2_4 = 11'B00000000000,
 _3I4274_$1I3863.CHAN_BOND_SEQ_2_USE = "FALSE",
 _3I4274_$1I3863.CHAN_BOND_SEQ_LEN = 1,
 _3I4274_$1I3863.CHAN_BOND_WAIT = 8,
 _3I4274_$1I3863.CLK_COR_INSERT_IDLE_FLAG = "FALSE",
 _3I4274_$1I3863.CLK_COR_KEEP_IDLE = TRUE,
 _3I4274_$1I3863.CLK_COR_REPEAT_WAIT = 0,
 _3I4274_$1I3863.CLK_COR_SEQ_1_1 = 00110111100,
 _3I4274_$1I3863.CLK_COR_SEQ_1_2 = 00011000101,
 _3I4274_$1I3863.CLK_COR_SEQ_1_3 = 11'B00000000000,
 _3I4274_$1I3863.CLK_COR_SEQ_1_4 = 11'B00000000000,
 _3I4274_$1I3863.CLK_COR_SEQ_2_1 = 00110111100,
 _3I4274_$1I3863.CLK_COR_SEQ_2_2 = 00001010000,
 _3I4274_$1I3863.CLK_COR_SEQ_2_3 = 11'B00000000000,
 _3I4274_$1I3863.CLK_COR_SEQ_2_4 = 11'B00000000000,
 _3I4274_$1I3863.CLK_COR_SEQ_2_USE = TRUE,
 _3I4274_$1I3863.CLK_COR_SEQ_LEN = 2,
 _3I4274_$1I3863.CLK_CORRECT_USE = "TRUE",
 _3I4274_$1I3863.COMMA_10B_MASK = 10'B1111111000,
 _3I4274_$1I3863.CRC_END_OF_PKT = "K29_7",
 _3I4274_$1I3863.CRC_FORMAT = "USER_MODE",
 _3I4274_$1I3863.CRC_START_OF_PKT = "K27_7",
 _3I4274_$1I3863.DEC_MCOMMA_DETECT = "TRUE",
 _3I4274_$1I3863.DEC_PCOMMA_DETECT = "TRUE",
 _3I4274_$1I3863.DEC_VALID_COMMA_ONLY = "TRUE",
 _3I4274_$1I3863.MCOMMA_10B_VALUE = 10'B1100000000,
 _3I4274_$1I3863.MCOMMA_DETECT = "TRUE",
 _3I4274_$1I3863.PCOMMA_10B_VALUE = 10'B0011111000,
 _3I4274_$1I3863.PCOMMA_DETECT = "TRUE",
 _3I4274_$1I3863.REF_CLK_V_SEL = 1,
 _3I4274_$1I3863.RX_BUFFER_USE = "TRUE",
 _3I4274_$1I3863.RX_CRC_USE = "FALSE",
 _3I4274_$1I3863.RX_DATA_WIDTH = 2,
 _3I4274_$1I3863.RX_DECODE_USE = "TRUE",
 _3I4274_$1I3863.RX_LOS_INVALID_INCR = 2,
 _3I4274_$1I3863.RX_LOS_THRESHOLD = 8,
 _3I4274_$1I3863.RX_LOSS_OF_SYNC_FSM = "TRUE",
 _3I4274_$1I3863.SERDES_10B = "FALSE",
 _3I4274_$1I3863.TERMINATION_IMP = 50,
 _3I4274_$1I3863.TX_BUFFER_USE = "TRUE",
 _3I4274_$1I3863.TX_CRC_FORCE_VALUE = 8'B11010110,
 _3I4274_$1I3863.TX_CRC_USE = "FALSE",
 _3I4274_$1I3863.TX_DATA_WIDTH = 2,
 _3I4274_$1I3863.TX_DIFF_CTRL = 400,
 _3I4274_$1I3863.TX_PREEMPHASIS = 0,
 _3I4243_$1I3863.ALIGN_COMMA_MSB = TRUE,
 _3I4243_$1I3863.CHAN_BOND_LIMIT = 16,
 _3I4243_$1I3863.CHAN_BOND_MODE = "OFF",
 _3I4243_$1I3863.CHAN_BOND_OFFSET = 8,
 _3I4243_$1I3863.CHAN_BOND_ONE_SHOT = "FALSE",
 _3I4243_$1I3863.CHAN_BOND_SEQ_1_1 = 11'B00000000000,
 _3I4243_$1I3863.CHAN_BOND_SEQ_1_2 = 11'B00000000000,
 _3I4243_$1I3863.CHAN_BOND_SEQ_1_3 = 11'B00000000000,
 _3I4243_$1I3863.CHAN_BOND_SEQ_1_4 = 11'B00000000000,
 _3I4243_$1I3863.CHAN_BOND_SEQ_2_1 = 11'B00000000000,
 _3I4243_$1I3863.CHAN_BOND_SEQ_2_2 = 11'B00000000000,
 _3I4243_$1I3863.CHAN_BOND_SEQ_2_3 = 11'B00000000000,
 _3I4243_$1I3863.CHAN_BOND_SEQ_2_4 = 11'B00000000000,
 _3I4243_$1I3863.CHAN_BOND_SEQ_2_USE = "FALSE",
 _3I4243_$1I3863.CHAN_BOND_SEQ_LEN = 1,
 _3I4243_$1I3863.CHAN_BOND_WAIT = 8,
 _3I4243_$1I3863.CLK_COR_INSERT_IDLE_FLAG = "FALSE",
 _3I4243_$1I3863.CLK_COR_KEEP_IDLE = TRUE,
 _3I4243_$1I3863.CLK_COR_REPEAT_WAIT = 0,
 _3I4243_$1I3863.CLK_COR_SEQ_1_1 = 00110111100,
 _3I4243_$1I3863.CLK_COR_SEQ_1_2 = 00011000101,
 _3I4243_$1I3863.CLK_COR_SEQ_1_3 = 11'B00000000000,
 _3I4243_$1I3863.CLK_COR_SEQ_1_4 = 11'B00000000000,
 _3I4243_$1I3863.CLK_COR_SEQ_2_1 = 00110111100,
 _3I4243_$1I3863.CLK_COR_SEQ_2_2 = 00001010000,
 _3I4243_$1I3863.CLK_COR_SEQ_2_3 = 11'B00000000000,
 _3I4243_$1I3863.CLK_COR_SEQ_2_4 = 11'B00000000000,
 _3I4243_$1I3863.CLK_COR_SEQ_2_USE = TRUE,
 _3I4243_$1I3863.CLK_COR_SEQ_LEN = 2,
 _3I4243_$1I3863.CLK_CORRECT_USE = "TRUE",
 _3I4243_$1I3863.COMMA_10B_MASK = 10'B1111111000,
 _3I4243_$1I3863.CRC_END_OF_PKT = "K29_7",
 _3I4243_$1I3863.CRC_FORMAT = "USER_MODE",
 _3I4243_$1I3863.CRC_START_OF_PKT = "K27_7",
 _3I4243_$1I3863.DEC_MCOMMA_DETECT = "TRUE",
 _3I4243_$1I3863.DEC_PCOMMA_DETECT = "TRUE",
 _3I4243_$1I3863.DEC_VALID_COMMA_ONLY = "TRUE",
 _3I4243_$1I3863.MCOMMA_10B_VALUE = 10'B1100000000,
 _3I4243_$1I3863.MCOMMA_DETECT = "TRUE",
 _3I4243_$1I3863.PCOMMA_10B_VALUE = 10'B0011111000,
 _3I4243_$1I3863.PCOMMA_DETECT = "TRUE",
 _3I4243_$1I3863.REF_CLK_V_SEL = 1,
 _3I4243_$1I3863.RX_BUFFER_USE = "TRUE",
 _3I4243_$1I3863.RX_CRC_USE = "FALSE",
 _3I4243_$1I3863.RX_DATA_WIDTH = 2,
 _3I4243_$1I3863.RX_DECODE_USE = "TRUE",
 _3I4243_$1I3863.RX_LOS_INVALID_INCR = 2,
 _3I4243_$1I3863.RX_LOS_THRESHOLD = 8,
 _3I4243_$1I3863.RX_LOSS_OF_SYNC_FSM = "TRUE",
 _3I4243_$1I3863.SERDES_10B = "FALSE",
 _3I4243_$1I3863.TERMINATION_IMP = 50,
 _3I4243_$1I3863.TX_BUFFER_USE = "TRUE",
 _3I4243_$1I3863.TX_CRC_FORCE_VALUE = 8'B11010110,
 _3I4243_$1I3863.TX_CRC_USE = "FALSE",
 _3I4243_$1I3863.TX_DATA_WIDTH = 2,
 _3I4243_$1I3863.TX_DIFF_CTRL = 400,
 _3I4243_$1I3863.TX_PREEMPHASIS = 0,
 _3I4142_$1I3863.ALIGN_COMMA_MSB = TRUE,
 _3I4142_$1I3863.CHAN_BOND_LIMIT = 16,
 _3I4142_$1I3863.CHAN_BOND_MODE = "OFF",
 _3I4142_$1I3863.CHAN_BOND_OFFSET = 8,
 _3I4142_$1I3863.CHAN_BOND_ONE_SHOT = "FALSE",
 _3I4142_$1I3863.CHAN_BOND_SEQ_1_1 = 11'B00000000000,
 _3I4142_$1I3863.CHAN_BOND_SEQ_1_2 = 11'B00000000000,
 _3I4142_$1I3863.CHAN_BOND_SEQ_1_3 = 11'B00000000000,
 _3I4142_$1I3863.CHAN_BOND_SEQ_1_4 = 11'B00000000000,
 _3I4142_$1I3863.CHAN_BOND_SEQ_2_1 = 11'B00000000000,
 _3I4142_$1I3863.CHAN_BOND_SEQ_2_2 = 11'B00000000000,
 _3I4142_$1I3863.CHAN_BOND_SEQ_2_3 = 11'B00000000000,
 _3I4142_$1I3863.CHAN_BOND_SEQ_2_4 = 11'B00000000000,
 _3I4142_$1I3863.CHAN_BOND_SEQ_2_USE = "FALSE",
 _3I4142_$1I3863.CHAN_BOND_SEQ_LEN = 1,
 _3I4142_$1I3863.CHAN_BOND_WAIT = 8,
 _3I4142_$1I3863.CLK_COR_INSERT_IDLE_FLAG = "FALSE",
 _3I4142_$1I3863.CLK_COR_KEEP_IDLE = TRUE,
 _3I4142_$1I3863.CLK_COR_REPEAT_WAIT = 0,
 _3I4142_$1I3863.CLK_COR_SEQ_1_1 = 00110111100,
 _3I4142_$1I3863.CLK_COR_SEQ_1_2 = 00011000101,
 _3I4142_$1I3863.CLK_COR_SEQ_1_3 = 11'B00000000000,
 _3I4142_$1I3863.CLK_COR_SEQ_1_4 = 11'B00000000000,
 _3I4142_$1I3863.CLK_COR_SEQ_2_1 = 00110111100,
 _3I4142_$1I3863.CLK_COR_SEQ_2_2 = 00001010000,
 _3I4142_$1I3863.CLK_COR_SEQ_2_3 = 11'B00000000000,
 _3I4142_$1I3863.CLK_COR_SEQ_2_4 = 11'B00000000000,
 _3I4142_$1I3863.CLK_COR_SEQ_2_USE = TRUE,
 _3I4142_$1I3863.CLK_COR_SEQ_LEN = 2,
 _3I4142_$1I3863.CLK_CORRECT_USE = "TRUE",
 _3I4142_$1I3863.COMMA_10B_MASK = 10'B1111111000,
 _3I4142_$1I3863.CRC_END_OF_PKT = "K29_7",
 _3I4142_$1I3863.CRC_FORMAT = "USER_MODE",
 _3I4142_$1I3863.CRC_START_OF_PKT = "K27_7",
 _3I4142_$1I3863.DEC_MCOMMA_DETECT = "TRUE",
 _3I4142_$1I3863.DEC_PCOMMA_DETECT = "TRUE",
 _3I4142_$1I3863.DEC_VALID_COMMA_ONLY = "TRUE",
 _3I4142_$1I3863.MCOMMA_10B_VALUE = 10'B1100000000,
 _3I4142_$1I3863.MCOMMA_DETECT = "TRUE",
 _3I4142_$1I3863.PCOMMA_10B_VALUE = 10'B0011111000,
 _3I4142_$1I3863.PCOMMA_DETECT = "TRUE",
 _3I4142_$1I3863.REF_CLK_V_SEL = 1,
 _3I4142_$1I3863.RX_BUFFER_USE = "TRUE",
 _3I4142_$1I3863.RX_CRC_USE = "FALSE",
 _3I4142_$1I3863.RX_DATA_WIDTH = 2,
 _3I4142_$1I3863.RX_DECODE_USE = "TRUE",
 _3I4142_$1I3863.RX_LOS_INVALID_INCR = 2,
 _3I4142_$1I3863.RX_LOS_THRESHOLD = 8,
 _3I4142_$1I3863.RX_LOSS_OF_SYNC_FSM = "TRUE",
 _3I4142_$1I3863.SERDES_10B = "FALSE",
 _3I4142_$1I3863.TERMINATION_IMP = 50,
 _3I4142_$1I3863.TX_BUFFER_USE = "TRUE",
 _3I4142_$1I3863.TX_CRC_FORCE_VALUE = 8'B11010110,
 _3I4142_$1I3863.TX_CRC_USE = "FALSE",
 _3I4142_$1I3863.TX_DATA_WIDTH = 2,
 _3I4142_$1I3863.TX_DIFF_CTRL = 400,
 _3I4142_$1I3863.TX_PREEMPHASIS = 0,
 _2I4609.CLK_FEEDBACK = "1X",
 _2I4609.CLKDV_DIVIDE = 2.0,
 _2I4609.CLKFX_DIVIDE = 1,
 _2I4609.CLKFX_MULTIPLY = 4,
 _2I4609.CLKIN_DIVIDE_BY_2 = "FALSE",
 _2I4609.CLKIN_PERIOD = 0.0,
 _2I4609.CLKOUT_PHASE_SHIFT = "NONE",
 _2I4609.DESKEW_ADJUST = "SYSTEM_SYNCHRONOUS",
 _2I4609.DFS_FREQUENCY_MODE = "LOW",
 _2I4609.DLL_FREQUENCY_MODE = "LOW",
 _2I4609.DSS_MODE = "NONE",
 _2I4609.DUTY_CYCLE_CORRECTION = "TRUE",
 _2I4609.FACTORY_JF = 16'HC080,
 _2I4609.PHASE_SHIFT = 0,
 _2I4609.STARTUP_WAIT = "FALSE",
 _2I4594.CLK_FEEDBACK = "1X",
 _2I4594.CLKDV_DIVIDE = 16.0,
 _2I4594.CLKFX_DIVIDE = 1,
 _2I4594.CLKFX_MULTIPLY = 4,
 _2I4594.CLKIN_DIVIDE_BY_2 = "FALSE",
 _2I4594.CLKIN_PERIOD = 0.0,
 _2I4594.CLKOUT_PHASE_SHIFT = "NONE",
 _2I4594.DESKEW_ADJUST = "SYSTEM_SYNCHRONOUS",
 _2I4594.DFS_FREQUENCY_MODE = "LOW",
 _2I4594.DLL_FREQUENCY_MODE = "LOW",
 _2I4594.DSS_MODE = "NONE",
 _2I4594.DUTY_CYCLE_CORRECTION = "TRUE",
 _2I4594.FACTORY_JF = 16'HC080,
 _2I4594.PHASE_SHIFT = 0,
 _2I4594.STARTUP_WAIT = TRUE,
 _1I4143_$1I4488_$1I4621.INIT_A = 9'H000,
 _1I4143_$1I4488_$1I4621.INIT_B = 18'H00000,
 _1I4143_$1I4488_$1I4621.SRVAL_A = 9'H000,
 _1I4143_$1I4488_$1I4621.SRVAL_B = 18'H00000,
 _1I4143_$1I4488_$1I4621.WRITE_MODE_A = "WRITE_FIRST",
 _1I4143_$1I4488_$1I4621.WRITE_MODE_B = "WRITE_FIRST",
 _1I4143_$1I4488_$1I4621.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4621.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_A = 9'H000,
 _1I4143_$1I4488_$1I4620.INIT_B = 18'H00000,
 _1I4143_$1I4488_$1I4620.SRVAL_A = 9'H000,
 _1I4143_$1I4488_$1I4620.SRVAL_B = 18'H00000,
 _1I4143_$1I4488_$1I4620.WRITE_MODE_A = "WRITE_FIRST",
 _1I4143_$1I4488_$1I4620.WRITE_MODE_B = "WRITE_FIRST",
 _1I4143_$1I4488_$1I4620.INIT_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_08 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_09 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_0A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_0B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_0C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_0D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_0E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_0F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_10 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_11 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_12 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_13 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_14 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_15 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_16 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_17 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_18 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_19 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_1A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_1B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_1C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_1D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_1E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_1F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_20 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_21 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_22 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_23 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_24 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_25 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_26 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_27 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_28 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_29 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_2A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_2B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_2C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_2D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_2E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_2F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_30 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_31 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_32 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_33 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_34 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_35 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_36 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_37 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_38 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_39 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_3A = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_3B = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_3C = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_3D = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_3E = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INIT_3F = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INITP_00 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INITP_01 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INITP_02 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INITP_03 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INITP_04 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INITP_05 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INITP_06 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4143_$1I4488_$1I4620.INITP_07 = 256'H0000000000000000000000000000000000000000000000000000000000000000,
 _1I4142_$1I3863.ALIGN_COMMA_MSB = TRUE,
 _1I4142_$1I3863.CHAN_BOND_LIMIT = 16,
 _1I4142_$1I3863.CHAN_BOND_MODE = "OFF",
 _1I4142_$1I3863.CHAN_BOND_OFFSET = 8,
 _1I4142_$1I3863.CHAN_BOND_ONE_SHOT = "FALSE",
 _1I4142_$1I3863.CHAN_BOND_SEQ_1_1 = 11'B00000000000,
 _1I4142_$1I3863.CHAN_BOND_SEQ_1_2 = 11'B00000000000,
 _1I4142_$1I3863.CHAN_BOND_SEQ_1_3 = 11'B00000000000,
 _1I4142_$1I3863.CHAN_BOND_SEQ_1_4 = 11'B00000000000,
 _1I4142_$1I3863.CHAN_BOND_SEQ_2_1 = 11'B00000000000,
 _1I4142_$1I3863.CHAN_BOND_SEQ_2_2 = 11'B00000000000,
 _1I4142_$1I3863.CHAN_BOND_SEQ_2_3 = 11'B00000000000,
 _1I4142_$1I3863.CHAN_BOND_SEQ_2_4 = 11'B00000000000,
 _1I4142_$1I3863.CHAN_BOND_SEQ_2_USE = "FALSE",
 _1I4142_$1I3863.CHAN_BOND_SEQ_LEN = 1,
 _1I4142_$1I3863.CHAN_BOND_WAIT = 8,
 _1I4142_$1I3863.CLK_COR_INSERT_IDLE_FLAG = "FALSE",
 _1I4142_$1I3863.CLK_COR_KEEP_IDLE = TRUE,
 _1I4142_$1I3863.CLK_COR_REPEAT_WAIT = 0,
 _1I4142_$1I3863.CLK_COR_SEQ_1_1 = 00110111100,
 _1I4142_$1I3863.CLK_COR_SEQ_1_2 = 00011000101,
 _1I4142_$1I3863.CLK_COR_SEQ_1_3 = 11'B00000000000,
 _1I4142_$1I3863.CLK_COR_SEQ_1_4 = 11'B00000000000,
 _1I4142_$1I3863.CLK_COR_SEQ_2_1 = 00110111100,
 _1I4142_$1I3863.CLK_COR_SEQ_2_2 = 00001010000,
 _1I4142_$1I3863.CLK_COR_SEQ_2_3 = 11'B00000000000,
 _1I4142_$1I3863.CLK_COR_SEQ_2_4 = 11'B00000000000,
 _1I4142_$1I3863.CLK_COR_SEQ_2_USE = TRUE,
 _1I4142_$1I3863.CLK_COR_SEQ_LEN = 2,
 _1I4142_$1I3863.CLK_CORRECT_USE = "TRUE",
 _1I4142_$1I3863.COMMA_10B_MASK = 10'B1111111000,
 _1I4142_$1I3863.CRC_END_OF_PKT = "K29_7",
 _1I4142_$1I3863.CRC_FORMAT = "USER_MODE",
 _1I4142_$1I3863.CRC_START_OF_PKT = "K27_7",
 _1I4142_$1I3863.DEC_MCOMMA_DETECT = "TRUE",
 _1I4142_$1I3863.DEC_PCOMMA_DETECT = "TRUE",
 _1I4142_$1I3863.DEC_VALID_COMMA_ONLY = "TRUE",
 _1I4142_$1I3863.MCOMMA_10B_VALUE = 10'B1100000000,
 _1I4142_$1I3863.MCOMMA_DETECT = "TRUE",
 _1I4142_$1I3863.PCOMMA_10B_VALUE = 10'B0011111000,
 _1I4142_$1I3863.PCOMMA_DETECT = "TRUE",
 _1I4142_$1I3863.REF_CLK_V_SEL = 1,
 _1I4142_$1I3863.RX_BUFFER_USE = "TRUE",
 _1I4142_$1I3863.RX_CRC_USE = "FALSE",
 _1I4142_$1I3863.RX_DATA_WIDTH = 2,
 _1I4142_$1I3863.RX_DECODE_USE = "TRUE",
 _1I4142_$1I3863.RX_LOS_INVALID_INCR = 2,
 _1I4142_$1I3863.RX_LOS_THRESHOLD = 8,
 _1I4142_$1I3863.RX_LOSS_OF_SYNC_FSM = "TRUE",
 _1I4142_$1I3863.SERDES_10B = "FALSE",
 _1I4142_$1I3863.TERMINATION_IMP = 50,
 _1I4142_$1I3863.TX_BUFFER_USE = "TRUE",
 _1I4142_$1I3863.TX_CRC_FORCE_VALUE = 8'B11010110,
 _1I4142_$1I3863.TX_CRC_USE = "FALSE",
 _1I4142_$1I3863.TX_DATA_WIDTH = 2,
 _1I4142_$1I3863.TX_DIFF_CTRL = 400,
 _1I4142_$1I3863.TX_PREEMPHASIS = 0;

 wire [7:0] _7I5013_$1I4488_$1I4621_DOA;

 wire [15:0] _7I5013_$1I4488_$1I4621_DOB;

 wire [0:0] _7I5013_$1I4488_$1I4621_DOPA;

 wire [1:0] _7I5013_$1I4488_$1I4621_DOPB;

 wire [10:0] _7I5013_$1I4488_$1I4621_ADDRA;
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1_10 (_7I5013_$1I4488_$1I4621_ADDRA[10], _7I5013_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1_9 (_7I5013_$1I4488_$1I4621_ADDRA[9], _7I5013_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1_8 (_7I5013_$1I4488_$1I4621_ADDRA[8], _7I5013_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1_7 (_7I5013_$1I4488_$1I4621_ADDRA[7], _7I5013_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1_6 (_7I5013_$1I4488_$1I4621_ADDRA[6], _7I5013_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1_5 (_7I5013_$1I4488_$1I4621_ADDRA[5], _7I5013_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1_4 (_7I5013_$1I4488_$1I4621_ADDRA[4], _7I5013_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1_3 (_7I5013_$1I4488_$1I4621_ADDRA[3], _7I5013_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1_2 (_7I5013_$1I4488_$1I4621_ADDRA[2], _7I5013_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1_1 (_7I5013_$1I4488_$1I4621_ADDRA[1], _7I5013_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1_0 (_7I5013_$1I4488_$1I4621_ADDRA[0], _7I5013_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _7I5013_$1I4488_$1I4621_ADDRB;
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_2_9 (_7I5013_$1I4488_$1I4621_ADDRB[9], _7I5013_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_2_8 (_7I5013_$1I4488_$1I4621_ADDRB[8], _7I5013_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_2_7 (_7I5013_$1I4488_$1I4621_ADDRB[7], _7I5013_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_2_6 (_7I5013_$1I4488_$1I4621_ADDRB[6], _7I5013_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_2_5 (_7I5013_$1I4488_$1I4621_ADDRB[5], _7I5013_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_2_4 (_7I5013_$1I4488_$1I4621_ADDRB[4], _7I5013_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_2_3 (_7I5013_$1I4488_$1I4621_ADDRB[3], _7I5013_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_2_2 (_7I5013_$1I4488_$1I4621_ADDRB[2], _7I5013_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_2_1 (_7I5013_$1I4488_$1I4621_ADDRB[1], _7I5013_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_2_0 (_7I5013_$1I4488_$1I4621_ADDRB[0], _7I5013_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _7I5013_$1I4488_$1I4621_CLKA;
 reg [1:16] _7I5013_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_3 (_7I5013_$1I4488_$1I4621_CLKA, _7I5013_$1I4488_$1I4621_CLKA__vlIN);

 wire  _7I5013_$1I4488_$1I4621_CLKB;
 reg [1:16] _7I5013_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_4 (_7I5013_$1I4488_$1I4621_CLKB, _7I5013_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _7I5013_$1I4488_$1I4621_DIA;
 reg [1:16] _7I5013_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_5_7 (_7I5013_$1I4488_$1I4621_DIA[7], _7I5013_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_5_6 (_7I5013_$1I4488_$1I4621_DIA[6], _7I5013_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_5_5 (_7I5013_$1I4488_$1I4621_DIA[5], _7I5013_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_5_4 (_7I5013_$1I4488_$1I4621_DIA[4], _7I5013_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_5_3 (_7I5013_$1I4488_$1I4621_DIA[3], _7I5013_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_5_2 (_7I5013_$1I4488_$1I4621_DIA[2], _7I5013_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_5_1 (_7I5013_$1I4488_$1I4621_DIA[1], _7I5013_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_5_0 (_7I5013_$1I4488_$1I4621_DIA[0], _7I5013_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _7I5013_$1I4488_$1I4621_DIB;
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_6_15 (_7I5013_$1I4488_$1I4621_DIB[15], _7I5013_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_6_14 (_7I5013_$1I4488_$1I4621_DIB[14], _7I5013_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_6_13 (_7I5013_$1I4488_$1I4621_DIB[13], _7I5013_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_6_12 (_7I5013_$1I4488_$1I4621_DIB[12], _7I5013_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_6_11 (_7I5013_$1I4488_$1I4621_DIB[11], _7I5013_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_6_10 (_7I5013_$1I4488_$1I4621_DIB[10], _7I5013_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_6_9 (_7I5013_$1I4488_$1I4621_DIB[9], _7I5013_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_6_8 (_7I5013_$1I4488_$1I4621_DIB[8], _7I5013_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_6_7 (_7I5013_$1I4488_$1I4621_DIB[7], _7I5013_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_6_6 (_7I5013_$1I4488_$1I4621_DIB[6], _7I5013_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_6_5 (_7I5013_$1I4488_$1I4621_DIB[5], _7I5013_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_6_4 (_7I5013_$1I4488_$1I4621_DIB[4], _7I5013_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_6_3 (_7I5013_$1I4488_$1I4621_DIB[3], _7I5013_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_6_2 (_7I5013_$1I4488_$1I4621_DIB[2], _7I5013_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_6_1 (_7I5013_$1I4488_$1I4621_DIB[1], _7I5013_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_6_0 (_7I5013_$1I4488_$1I4621_DIB[0], _7I5013_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _7I5013_$1I4488_$1I4621_DIPA;
 reg [1:16] _7I5013_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_7_0 (_7I5013_$1I4488_$1I4621_DIPA[0], _7I5013_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _7I5013_$1I4488_$1I4621_DIPB;
 reg [1:16] _7I5013_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_8_1 (_7I5013_$1I4488_$1I4621_DIPB[1], _7I5013_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_8_0 (_7I5013_$1I4488_$1I4621_DIPB[0], _7I5013_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _7I5013_$1I4488_$1I4621_ENA;
 reg [1:16] _7I5013_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_9 (_7I5013_$1I4488_$1I4621_ENA, _7I5013_$1I4488_$1I4621_ENA__vlIN);

 wire  _7I5013_$1I4488_$1I4621_ENB;
 reg [1:16] _7I5013_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_10 (_7I5013_$1I4488_$1I4621_ENB, _7I5013_$1I4488_$1I4621_ENB__vlIN);

 wire  _7I5013_$1I4488_$1I4621_SSRA;
 reg [1:16] _7I5013_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_11 (_7I5013_$1I4488_$1I4621_SSRA, _7I5013_$1I4488_$1I4621_SSRA__vlIN);

 wire  _7I5013_$1I4488_$1I4621_SSRB;
 reg [1:16] _7I5013_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_12 (_7I5013_$1I4488_$1I4621_SSRB, _7I5013_$1I4488_$1I4621_SSRB__vlIN);

 wire  _7I5013_$1I4488_$1I4621_WEA;
 reg [1:16] _7I5013_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_13 (_7I5013_$1I4488_$1I4621_WEA, _7I5013_$1I4488_$1I4621_WEA__vlIN);

 wire  _7I5013_$1I4488_$1I4621_WEB;
 reg [1:16] _7I5013_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_14 (_7I5013_$1I4488_$1I4621_WEB, _7I5013_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _7I5013_$1I4488_$1I4621 ( _7I5013_$1I4488_$1I4621_DOA , _7I5013_$1I4488_$1I4621_DOB , _7I5013_$1I4488_$1I4621_DOPA , _7I5013_$1I4488_$1I4621_DOPB , _7I5013_$1I4488_$1I4621_ADDRA , _7I5013_$1I4488_$1I4621_ADDRB , _7I5013_$1I4488_$1I4621_CLKA , _7I5013_$1I4488_$1I4621_CLKB , _7I5013_$1I4488_$1I4621_DIA , _7I5013_$1I4488_$1I4621_DIB , _7I5013_$1I4488_$1I4621_DIPA , _7I5013_$1I4488_$1I4621_DIPB , _7I5013_$1I4488_$1I4621_ENA , _7I5013_$1I4488_$1I4621_ENB , _7I5013_$1I4488_$1I4621_SSRA , _7I5013_$1I4488_$1I4621_SSRB , _7I5013_$1I4488_$1I4621_WEA , _7I5013_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _7I5013_$1I4488_$1I4620_DOA;

 wire [15:0] _7I5013_$1I4488_$1I4620_DOB;

 wire [0:0] _7I5013_$1I4488_$1I4620_DOPA;

 wire [1:0] _7I5013_$1I4488_$1I4620_DOPB;

 wire [10:0] _7I5013_$1I4488_$1I4620_ADDRA;
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_15_10 (_7I5013_$1I4488_$1I4620_ADDRA[10], _7I5013_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_15_9 (_7I5013_$1I4488_$1I4620_ADDRA[9], _7I5013_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_15_8 (_7I5013_$1I4488_$1I4620_ADDRA[8], _7I5013_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_15_7 (_7I5013_$1I4488_$1I4620_ADDRA[7], _7I5013_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_15_6 (_7I5013_$1I4488_$1I4620_ADDRA[6], _7I5013_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_15_5 (_7I5013_$1I4488_$1I4620_ADDRA[5], _7I5013_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_15_4 (_7I5013_$1I4488_$1I4620_ADDRA[4], _7I5013_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_15_3 (_7I5013_$1I4488_$1I4620_ADDRA[3], _7I5013_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_15_2 (_7I5013_$1I4488_$1I4620_ADDRA[2], _7I5013_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_15_1 (_7I5013_$1I4488_$1I4620_ADDRA[1], _7I5013_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_15_0 (_7I5013_$1I4488_$1I4620_ADDRA[0], _7I5013_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _7I5013_$1I4488_$1I4620_ADDRB;
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_16_9 (_7I5013_$1I4488_$1I4620_ADDRB[9], _7I5013_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_16_8 (_7I5013_$1I4488_$1I4620_ADDRB[8], _7I5013_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_16_7 (_7I5013_$1I4488_$1I4620_ADDRB[7], _7I5013_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_16_6 (_7I5013_$1I4488_$1I4620_ADDRB[6], _7I5013_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_16_5 (_7I5013_$1I4488_$1I4620_ADDRB[5], _7I5013_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_16_4 (_7I5013_$1I4488_$1I4620_ADDRB[4], _7I5013_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_16_3 (_7I5013_$1I4488_$1I4620_ADDRB[3], _7I5013_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_16_2 (_7I5013_$1I4488_$1I4620_ADDRB[2], _7I5013_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_16_1 (_7I5013_$1I4488_$1I4620_ADDRB[1], _7I5013_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_16_0 (_7I5013_$1I4488_$1I4620_ADDRB[0], _7I5013_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _7I5013_$1I4488_$1I4620_CLKA;
 reg [1:16] _7I5013_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_17 (_7I5013_$1I4488_$1I4620_CLKA, _7I5013_$1I4488_$1I4620_CLKA__vlIN);

 wire  _7I5013_$1I4488_$1I4620_CLKB;
 reg [1:16] _7I5013_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_18 (_7I5013_$1I4488_$1I4620_CLKB, _7I5013_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _7I5013_$1I4488_$1I4620_DIA;
 reg [1:16] _7I5013_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_19_7 (_7I5013_$1I4488_$1I4620_DIA[7], _7I5013_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_19_6 (_7I5013_$1I4488_$1I4620_DIA[6], _7I5013_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_19_5 (_7I5013_$1I4488_$1I4620_DIA[5], _7I5013_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_19_4 (_7I5013_$1I4488_$1I4620_DIA[4], _7I5013_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_19_3 (_7I5013_$1I4488_$1I4620_DIA[3], _7I5013_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_19_2 (_7I5013_$1I4488_$1I4620_DIA[2], _7I5013_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_19_1 (_7I5013_$1I4488_$1I4620_DIA[1], _7I5013_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_19_0 (_7I5013_$1I4488_$1I4620_DIA[0], _7I5013_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _7I5013_$1I4488_$1I4620_DIB;
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_20_15 (_7I5013_$1I4488_$1I4620_DIB[15], _7I5013_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_20_14 (_7I5013_$1I4488_$1I4620_DIB[14], _7I5013_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_20_13 (_7I5013_$1I4488_$1I4620_DIB[13], _7I5013_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_20_12 (_7I5013_$1I4488_$1I4620_DIB[12], _7I5013_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_20_11 (_7I5013_$1I4488_$1I4620_DIB[11], _7I5013_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_20_10 (_7I5013_$1I4488_$1I4620_DIB[10], _7I5013_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_20_9 (_7I5013_$1I4488_$1I4620_DIB[9], _7I5013_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_20_8 (_7I5013_$1I4488_$1I4620_DIB[8], _7I5013_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_20_7 (_7I5013_$1I4488_$1I4620_DIB[7], _7I5013_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_20_6 (_7I5013_$1I4488_$1I4620_DIB[6], _7I5013_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_20_5 (_7I5013_$1I4488_$1I4620_DIB[5], _7I5013_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_20_4 (_7I5013_$1I4488_$1I4620_DIB[4], _7I5013_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_20_3 (_7I5013_$1I4488_$1I4620_DIB[3], _7I5013_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_20_2 (_7I5013_$1I4488_$1I4620_DIB[2], _7I5013_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_20_1 (_7I5013_$1I4488_$1I4620_DIB[1], _7I5013_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_20_0 (_7I5013_$1I4488_$1I4620_DIB[0], _7I5013_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _7I5013_$1I4488_$1I4620_DIPA;
 reg [1:16] _7I5013_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_21_0 (_7I5013_$1I4488_$1I4620_DIPA[0], _7I5013_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _7I5013_$1I4488_$1I4620_DIPB;
 reg [1:16] _7I5013_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_22_1 (_7I5013_$1I4488_$1I4620_DIPB[1], _7I5013_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _7I5013_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_22_0 (_7I5013_$1I4488_$1I4620_DIPB[0], _7I5013_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _7I5013_$1I4488_$1I4620_ENA;
 reg [1:16] _7I5013_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_23 (_7I5013_$1I4488_$1I4620_ENA, _7I5013_$1I4488_$1I4620_ENA__vlIN);

 wire  _7I5013_$1I4488_$1I4620_ENB;
 reg [1:16] _7I5013_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_24 (_7I5013_$1I4488_$1I4620_ENB, _7I5013_$1I4488_$1I4620_ENB__vlIN);

 wire  _7I5013_$1I4488_$1I4620_SSRA;
 reg [1:16] _7I5013_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_25 (_7I5013_$1I4488_$1I4620_SSRA, _7I5013_$1I4488_$1I4620_SSRA__vlIN);

 wire  _7I5013_$1I4488_$1I4620_SSRB;
 reg [1:16] _7I5013_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_26 (_7I5013_$1I4488_$1I4620_SSRB, _7I5013_$1I4488_$1I4620_SSRB__vlIN);

 wire  _7I5013_$1I4488_$1I4620_WEA;
 reg [1:16] _7I5013_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_27 (_7I5013_$1I4488_$1I4620_WEA, _7I5013_$1I4488_$1I4620_WEA__vlIN);

 wire  _7I5013_$1I4488_$1I4620_WEB;
 reg [1:16] _7I5013_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_28 (_7I5013_$1I4488_$1I4620_WEB, _7I5013_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _7I5013_$1I4488_$1I4620 ( _7I5013_$1I4488_$1I4620_DOA , _7I5013_$1I4488_$1I4620_DOB , _7I5013_$1I4488_$1I4620_DOPA , _7I5013_$1I4488_$1I4620_DOPB , _7I5013_$1I4488_$1I4620_ADDRA , _7I5013_$1I4488_$1I4620_ADDRB , _7I5013_$1I4488_$1I4620_CLKA , _7I5013_$1I4488_$1I4620_CLKB , _7I5013_$1I4488_$1I4620_DIA , _7I5013_$1I4488_$1I4620_DIB , _7I5013_$1I4488_$1I4620_DIPA , _7I5013_$1I4488_$1I4620_DIPB , _7I5013_$1I4488_$1I4620_ENA , _7I5013_$1I4488_$1I4620_ENB , _7I5013_$1I4488_$1I4620_SSRA , _7I5013_$1I4488_$1I4620_SSRB , _7I5013_$1I4488_$1I4620_WEA , _7I5013_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4974_$1I4488_$1I4621_DOA;

 wire [15:0] _7I4974_$1I4488_$1I4621_DOB;

 wire [0:0] _7I4974_$1I4488_$1I4621_DOPA;

 wire [1:0] _7I4974_$1I4488_$1I4621_DOPB;

 wire [10:0] _7I4974_$1I4488_$1I4621_ADDRA;
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_29_10 (_7I4974_$1I4488_$1I4621_ADDRA[10], _7I4974_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_29_9 (_7I4974_$1I4488_$1I4621_ADDRA[9], _7I4974_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_29_8 (_7I4974_$1I4488_$1I4621_ADDRA[8], _7I4974_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_29_7 (_7I4974_$1I4488_$1I4621_ADDRA[7], _7I4974_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_29_6 (_7I4974_$1I4488_$1I4621_ADDRA[6], _7I4974_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_29_5 (_7I4974_$1I4488_$1I4621_ADDRA[5], _7I4974_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_29_4 (_7I4974_$1I4488_$1I4621_ADDRA[4], _7I4974_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_29_3 (_7I4974_$1I4488_$1I4621_ADDRA[3], _7I4974_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_29_2 (_7I4974_$1I4488_$1I4621_ADDRA[2], _7I4974_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_29_1 (_7I4974_$1I4488_$1I4621_ADDRA[1], _7I4974_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_29_0 (_7I4974_$1I4488_$1I4621_ADDRA[0], _7I4974_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _7I4974_$1I4488_$1I4621_ADDRB;
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_30_9 (_7I4974_$1I4488_$1I4621_ADDRB[9], _7I4974_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_30_8 (_7I4974_$1I4488_$1I4621_ADDRB[8], _7I4974_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_30_7 (_7I4974_$1I4488_$1I4621_ADDRB[7], _7I4974_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_30_6 (_7I4974_$1I4488_$1I4621_ADDRB[6], _7I4974_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_30_5 (_7I4974_$1I4488_$1I4621_ADDRB[5], _7I4974_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_30_4 (_7I4974_$1I4488_$1I4621_ADDRB[4], _7I4974_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_30_3 (_7I4974_$1I4488_$1I4621_ADDRB[3], _7I4974_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_30_2 (_7I4974_$1I4488_$1I4621_ADDRB[2], _7I4974_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_30_1 (_7I4974_$1I4488_$1I4621_ADDRB[1], _7I4974_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_30_0 (_7I4974_$1I4488_$1I4621_ADDRB[0], _7I4974_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _7I4974_$1I4488_$1I4621_CLKA;
 reg [1:16] _7I4974_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_31 (_7I4974_$1I4488_$1I4621_CLKA, _7I4974_$1I4488_$1I4621_CLKA__vlIN);

 wire  _7I4974_$1I4488_$1I4621_CLKB;
 reg [1:16] _7I4974_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_32 (_7I4974_$1I4488_$1I4621_CLKB, _7I4974_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _7I4974_$1I4488_$1I4621_DIA;
 reg [1:16] _7I4974_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_33_7 (_7I4974_$1I4488_$1I4621_DIA[7], _7I4974_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_33_6 (_7I4974_$1I4488_$1I4621_DIA[6], _7I4974_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_33_5 (_7I4974_$1I4488_$1I4621_DIA[5], _7I4974_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_33_4 (_7I4974_$1I4488_$1I4621_DIA[4], _7I4974_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_33_3 (_7I4974_$1I4488_$1I4621_DIA[3], _7I4974_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_33_2 (_7I4974_$1I4488_$1I4621_DIA[2], _7I4974_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_33_1 (_7I4974_$1I4488_$1I4621_DIA[1], _7I4974_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_33_0 (_7I4974_$1I4488_$1I4621_DIA[0], _7I4974_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _7I4974_$1I4488_$1I4621_DIB;
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_34_15 (_7I4974_$1I4488_$1I4621_DIB[15], _7I4974_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_34_14 (_7I4974_$1I4488_$1I4621_DIB[14], _7I4974_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_34_13 (_7I4974_$1I4488_$1I4621_DIB[13], _7I4974_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_34_12 (_7I4974_$1I4488_$1I4621_DIB[12], _7I4974_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_34_11 (_7I4974_$1I4488_$1I4621_DIB[11], _7I4974_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_34_10 (_7I4974_$1I4488_$1I4621_DIB[10], _7I4974_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_34_9 (_7I4974_$1I4488_$1I4621_DIB[9], _7I4974_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_34_8 (_7I4974_$1I4488_$1I4621_DIB[8], _7I4974_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_34_7 (_7I4974_$1I4488_$1I4621_DIB[7], _7I4974_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_34_6 (_7I4974_$1I4488_$1I4621_DIB[6], _7I4974_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_34_5 (_7I4974_$1I4488_$1I4621_DIB[5], _7I4974_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_34_4 (_7I4974_$1I4488_$1I4621_DIB[4], _7I4974_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_34_3 (_7I4974_$1I4488_$1I4621_DIB[3], _7I4974_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_34_2 (_7I4974_$1I4488_$1I4621_DIB[2], _7I4974_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_34_1 (_7I4974_$1I4488_$1I4621_DIB[1], _7I4974_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_34_0 (_7I4974_$1I4488_$1I4621_DIB[0], _7I4974_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _7I4974_$1I4488_$1I4621_DIPA;
 reg [1:16] _7I4974_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_35_0 (_7I4974_$1I4488_$1I4621_DIPA[0], _7I4974_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _7I4974_$1I4488_$1I4621_DIPB;
 reg [1:16] _7I4974_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_36_1 (_7I4974_$1I4488_$1I4621_DIPB[1], _7I4974_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_36_0 (_7I4974_$1I4488_$1I4621_DIPB[0], _7I4974_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _7I4974_$1I4488_$1I4621_ENA;
 reg [1:16] _7I4974_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_37 (_7I4974_$1I4488_$1I4621_ENA, _7I4974_$1I4488_$1I4621_ENA__vlIN);

 wire  _7I4974_$1I4488_$1I4621_ENB;
 reg [1:16] _7I4974_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_38 (_7I4974_$1I4488_$1I4621_ENB, _7I4974_$1I4488_$1I4621_ENB__vlIN);

 wire  _7I4974_$1I4488_$1I4621_SSRA;
 reg [1:16] _7I4974_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_39 (_7I4974_$1I4488_$1I4621_SSRA, _7I4974_$1I4488_$1I4621_SSRA__vlIN);

 wire  _7I4974_$1I4488_$1I4621_SSRB;
 reg [1:16] _7I4974_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_40 (_7I4974_$1I4488_$1I4621_SSRB, _7I4974_$1I4488_$1I4621_SSRB__vlIN);

 wire  _7I4974_$1I4488_$1I4621_WEA;
 reg [1:16] _7I4974_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_41 (_7I4974_$1I4488_$1I4621_WEA, _7I4974_$1I4488_$1I4621_WEA__vlIN);

 wire  _7I4974_$1I4488_$1I4621_WEB;
 reg [1:16] _7I4974_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_42 (_7I4974_$1I4488_$1I4621_WEB, _7I4974_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _7I4974_$1I4488_$1I4621 ( _7I4974_$1I4488_$1I4621_DOA , _7I4974_$1I4488_$1I4621_DOB , _7I4974_$1I4488_$1I4621_DOPA , _7I4974_$1I4488_$1I4621_DOPB , _7I4974_$1I4488_$1I4621_ADDRA , _7I4974_$1I4488_$1I4621_ADDRB , _7I4974_$1I4488_$1I4621_CLKA , _7I4974_$1I4488_$1I4621_CLKB , _7I4974_$1I4488_$1I4621_DIA , _7I4974_$1I4488_$1I4621_DIB , _7I4974_$1I4488_$1I4621_DIPA , _7I4974_$1I4488_$1I4621_DIPB , _7I4974_$1I4488_$1I4621_ENA , _7I4974_$1I4488_$1I4621_ENB , _7I4974_$1I4488_$1I4621_SSRA , _7I4974_$1I4488_$1I4621_SSRB , _7I4974_$1I4488_$1I4621_WEA , _7I4974_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4974_$1I4488_$1I4620_DOA;

 wire [15:0] _7I4974_$1I4488_$1I4620_DOB;

 wire [0:0] _7I4974_$1I4488_$1I4620_DOPA;

 wire [1:0] _7I4974_$1I4488_$1I4620_DOPB;

 wire [10:0] _7I4974_$1I4488_$1I4620_ADDRA;
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_43_10 (_7I4974_$1I4488_$1I4620_ADDRA[10], _7I4974_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_43_9 (_7I4974_$1I4488_$1I4620_ADDRA[9], _7I4974_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_43_8 (_7I4974_$1I4488_$1I4620_ADDRA[8], _7I4974_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_43_7 (_7I4974_$1I4488_$1I4620_ADDRA[7], _7I4974_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_43_6 (_7I4974_$1I4488_$1I4620_ADDRA[6], _7I4974_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_43_5 (_7I4974_$1I4488_$1I4620_ADDRA[5], _7I4974_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_43_4 (_7I4974_$1I4488_$1I4620_ADDRA[4], _7I4974_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_43_3 (_7I4974_$1I4488_$1I4620_ADDRA[3], _7I4974_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_43_2 (_7I4974_$1I4488_$1I4620_ADDRA[2], _7I4974_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_43_1 (_7I4974_$1I4488_$1I4620_ADDRA[1], _7I4974_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_43_0 (_7I4974_$1I4488_$1I4620_ADDRA[0], _7I4974_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _7I4974_$1I4488_$1I4620_ADDRB;
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_44_9 (_7I4974_$1I4488_$1I4620_ADDRB[9], _7I4974_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_44_8 (_7I4974_$1I4488_$1I4620_ADDRB[8], _7I4974_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_44_7 (_7I4974_$1I4488_$1I4620_ADDRB[7], _7I4974_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_44_6 (_7I4974_$1I4488_$1I4620_ADDRB[6], _7I4974_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_44_5 (_7I4974_$1I4488_$1I4620_ADDRB[5], _7I4974_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_44_4 (_7I4974_$1I4488_$1I4620_ADDRB[4], _7I4974_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_44_3 (_7I4974_$1I4488_$1I4620_ADDRB[3], _7I4974_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_44_2 (_7I4974_$1I4488_$1I4620_ADDRB[2], _7I4974_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_44_1 (_7I4974_$1I4488_$1I4620_ADDRB[1], _7I4974_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_44_0 (_7I4974_$1I4488_$1I4620_ADDRB[0], _7I4974_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _7I4974_$1I4488_$1I4620_CLKA;
 reg [1:16] _7I4974_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_45 (_7I4974_$1I4488_$1I4620_CLKA, _7I4974_$1I4488_$1I4620_CLKA__vlIN);

 wire  _7I4974_$1I4488_$1I4620_CLKB;
 reg [1:16] _7I4974_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_46 (_7I4974_$1I4488_$1I4620_CLKB, _7I4974_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _7I4974_$1I4488_$1I4620_DIA;
 reg [1:16] _7I4974_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_47_7 (_7I4974_$1I4488_$1I4620_DIA[7], _7I4974_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_47_6 (_7I4974_$1I4488_$1I4620_DIA[6], _7I4974_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_47_5 (_7I4974_$1I4488_$1I4620_DIA[5], _7I4974_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_47_4 (_7I4974_$1I4488_$1I4620_DIA[4], _7I4974_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_47_3 (_7I4974_$1I4488_$1I4620_DIA[3], _7I4974_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_47_2 (_7I4974_$1I4488_$1I4620_DIA[2], _7I4974_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_47_1 (_7I4974_$1I4488_$1I4620_DIA[1], _7I4974_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_47_0 (_7I4974_$1I4488_$1I4620_DIA[0], _7I4974_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _7I4974_$1I4488_$1I4620_DIB;
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_48_15 (_7I4974_$1I4488_$1I4620_DIB[15], _7I4974_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_48_14 (_7I4974_$1I4488_$1I4620_DIB[14], _7I4974_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_48_13 (_7I4974_$1I4488_$1I4620_DIB[13], _7I4974_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_48_12 (_7I4974_$1I4488_$1I4620_DIB[12], _7I4974_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_48_11 (_7I4974_$1I4488_$1I4620_DIB[11], _7I4974_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_48_10 (_7I4974_$1I4488_$1I4620_DIB[10], _7I4974_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_48_9 (_7I4974_$1I4488_$1I4620_DIB[9], _7I4974_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_48_8 (_7I4974_$1I4488_$1I4620_DIB[8], _7I4974_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_48_7 (_7I4974_$1I4488_$1I4620_DIB[7], _7I4974_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_48_6 (_7I4974_$1I4488_$1I4620_DIB[6], _7I4974_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_48_5 (_7I4974_$1I4488_$1I4620_DIB[5], _7I4974_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_48_4 (_7I4974_$1I4488_$1I4620_DIB[4], _7I4974_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_48_3 (_7I4974_$1I4488_$1I4620_DIB[3], _7I4974_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_48_2 (_7I4974_$1I4488_$1I4620_DIB[2], _7I4974_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_48_1 (_7I4974_$1I4488_$1I4620_DIB[1], _7I4974_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_48_0 (_7I4974_$1I4488_$1I4620_DIB[0], _7I4974_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _7I4974_$1I4488_$1I4620_DIPA;
 reg [1:16] _7I4974_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_49_0 (_7I4974_$1I4488_$1I4620_DIPA[0], _7I4974_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _7I4974_$1I4488_$1I4620_DIPB;
 reg [1:16] _7I4974_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_50_1 (_7I4974_$1I4488_$1I4620_DIPB[1], _7I4974_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _7I4974_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_50_0 (_7I4974_$1I4488_$1I4620_DIPB[0], _7I4974_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _7I4974_$1I4488_$1I4620_ENA;
 reg [1:16] _7I4974_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_51 (_7I4974_$1I4488_$1I4620_ENA, _7I4974_$1I4488_$1I4620_ENA__vlIN);

 wire  _7I4974_$1I4488_$1I4620_ENB;
 reg [1:16] _7I4974_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_52 (_7I4974_$1I4488_$1I4620_ENB, _7I4974_$1I4488_$1I4620_ENB__vlIN);

 wire  _7I4974_$1I4488_$1I4620_SSRA;
 reg [1:16] _7I4974_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_53 (_7I4974_$1I4488_$1I4620_SSRA, _7I4974_$1I4488_$1I4620_SSRA__vlIN);

 wire  _7I4974_$1I4488_$1I4620_SSRB;
 reg [1:16] _7I4974_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_54 (_7I4974_$1I4488_$1I4620_SSRB, _7I4974_$1I4488_$1I4620_SSRB__vlIN);

 wire  _7I4974_$1I4488_$1I4620_WEA;
 reg [1:16] _7I4974_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_55 (_7I4974_$1I4488_$1I4620_WEA, _7I4974_$1I4488_$1I4620_WEA__vlIN);

 wire  _7I4974_$1I4488_$1I4620_WEB;
 reg [1:16] _7I4974_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_56 (_7I4974_$1I4488_$1I4620_WEB, _7I4974_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _7I4974_$1I4488_$1I4620 ( _7I4974_$1I4488_$1I4620_DOA , _7I4974_$1I4488_$1I4620_DOB , _7I4974_$1I4488_$1I4620_DOPA , _7I4974_$1I4488_$1I4620_DOPB , _7I4974_$1I4488_$1I4620_ADDRA , _7I4974_$1I4488_$1I4620_ADDRB , _7I4974_$1I4488_$1I4620_CLKA , _7I4974_$1I4488_$1I4620_CLKB , _7I4974_$1I4488_$1I4620_DIA , _7I4974_$1I4488_$1I4620_DIB , _7I4974_$1I4488_$1I4620_DIPA , _7I4974_$1I4488_$1I4620_DIPB , _7I4974_$1I4488_$1I4620_ENA , _7I4974_$1I4488_$1I4620_ENB , _7I4974_$1I4488_$1I4620_SSRA , _7I4974_$1I4488_$1I4620_SSRB , _7I4974_$1I4488_$1I4620_WEA , _7I4974_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4863_$1I4488_$1I4621_DOA;

 wire [15:0] _7I4863_$1I4488_$1I4621_DOB;

 wire [0:0] _7I4863_$1I4488_$1I4621_DOPA;

 wire [1:0] _7I4863_$1I4488_$1I4621_DOPB;

 wire [10:0] _7I4863_$1I4488_$1I4621_ADDRA;
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_57_10 (_7I4863_$1I4488_$1I4621_ADDRA[10], _7I4863_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_57_9 (_7I4863_$1I4488_$1I4621_ADDRA[9], _7I4863_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_57_8 (_7I4863_$1I4488_$1I4621_ADDRA[8], _7I4863_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_57_7 (_7I4863_$1I4488_$1I4621_ADDRA[7], _7I4863_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_57_6 (_7I4863_$1I4488_$1I4621_ADDRA[6], _7I4863_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_57_5 (_7I4863_$1I4488_$1I4621_ADDRA[5], _7I4863_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_57_4 (_7I4863_$1I4488_$1I4621_ADDRA[4], _7I4863_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_57_3 (_7I4863_$1I4488_$1I4621_ADDRA[3], _7I4863_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_57_2 (_7I4863_$1I4488_$1I4621_ADDRA[2], _7I4863_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_57_1 (_7I4863_$1I4488_$1I4621_ADDRA[1], _7I4863_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_57_0 (_7I4863_$1I4488_$1I4621_ADDRA[0], _7I4863_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _7I4863_$1I4488_$1I4621_ADDRB;
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_58_9 (_7I4863_$1I4488_$1I4621_ADDRB[9], _7I4863_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_58_8 (_7I4863_$1I4488_$1I4621_ADDRB[8], _7I4863_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_58_7 (_7I4863_$1I4488_$1I4621_ADDRB[7], _7I4863_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_58_6 (_7I4863_$1I4488_$1I4621_ADDRB[6], _7I4863_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_58_5 (_7I4863_$1I4488_$1I4621_ADDRB[5], _7I4863_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_58_4 (_7I4863_$1I4488_$1I4621_ADDRB[4], _7I4863_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_58_3 (_7I4863_$1I4488_$1I4621_ADDRB[3], _7I4863_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_58_2 (_7I4863_$1I4488_$1I4621_ADDRB[2], _7I4863_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_58_1 (_7I4863_$1I4488_$1I4621_ADDRB[1], _7I4863_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_58_0 (_7I4863_$1I4488_$1I4621_ADDRB[0], _7I4863_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _7I4863_$1I4488_$1I4621_CLKA;
 reg [1:16] _7I4863_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_59 (_7I4863_$1I4488_$1I4621_CLKA, _7I4863_$1I4488_$1I4621_CLKA__vlIN);

 wire  _7I4863_$1I4488_$1I4621_CLKB;
 reg [1:16] _7I4863_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_60 (_7I4863_$1I4488_$1I4621_CLKB, _7I4863_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _7I4863_$1I4488_$1I4621_DIA;
 reg [1:16] _7I4863_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_61_7 (_7I4863_$1I4488_$1I4621_DIA[7], _7I4863_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_61_6 (_7I4863_$1I4488_$1I4621_DIA[6], _7I4863_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_61_5 (_7I4863_$1I4488_$1I4621_DIA[5], _7I4863_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_61_4 (_7I4863_$1I4488_$1I4621_DIA[4], _7I4863_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_61_3 (_7I4863_$1I4488_$1I4621_DIA[3], _7I4863_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_61_2 (_7I4863_$1I4488_$1I4621_DIA[2], _7I4863_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_61_1 (_7I4863_$1I4488_$1I4621_DIA[1], _7I4863_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_61_0 (_7I4863_$1I4488_$1I4621_DIA[0], _7I4863_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _7I4863_$1I4488_$1I4621_DIB;
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_62_15 (_7I4863_$1I4488_$1I4621_DIB[15], _7I4863_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_62_14 (_7I4863_$1I4488_$1I4621_DIB[14], _7I4863_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_62_13 (_7I4863_$1I4488_$1I4621_DIB[13], _7I4863_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_62_12 (_7I4863_$1I4488_$1I4621_DIB[12], _7I4863_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_62_11 (_7I4863_$1I4488_$1I4621_DIB[11], _7I4863_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_62_10 (_7I4863_$1I4488_$1I4621_DIB[10], _7I4863_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_62_9 (_7I4863_$1I4488_$1I4621_DIB[9], _7I4863_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_62_8 (_7I4863_$1I4488_$1I4621_DIB[8], _7I4863_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_62_7 (_7I4863_$1I4488_$1I4621_DIB[7], _7I4863_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_62_6 (_7I4863_$1I4488_$1I4621_DIB[6], _7I4863_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_62_5 (_7I4863_$1I4488_$1I4621_DIB[5], _7I4863_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_62_4 (_7I4863_$1I4488_$1I4621_DIB[4], _7I4863_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_62_3 (_7I4863_$1I4488_$1I4621_DIB[3], _7I4863_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_62_2 (_7I4863_$1I4488_$1I4621_DIB[2], _7I4863_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_62_1 (_7I4863_$1I4488_$1I4621_DIB[1], _7I4863_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_62_0 (_7I4863_$1I4488_$1I4621_DIB[0], _7I4863_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _7I4863_$1I4488_$1I4621_DIPA;
 reg [1:16] _7I4863_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_63_0 (_7I4863_$1I4488_$1I4621_DIPA[0], _7I4863_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _7I4863_$1I4488_$1I4621_DIPB;
 reg [1:16] _7I4863_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_64_1 (_7I4863_$1I4488_$1I4621_DIPB[1], _7I4863_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_64_0 (_7I4863_$1I4488_$1I4621_DIPB[0], _7I4863_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _7I4863_$1I4488_$1I4621_ENA;
 reg [1:16] _7I4863_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_65 (_7I4863_$1I4488_$1I4621_ENA, _7I4863_$1I4488_$1I4621_ENA__vlIN);

 wire  _7I4863_$1I4488_$1I4621_ENB;
 reg [1:16] _7I4863_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_66 (_7I4863_$1I4488_$1I4621_ENB, _7I4863_$1I4488_$1I4621_ENB__vlIN);

 wire  _7I4863_$1I4488_$1I4621_SSRA;
 reg [1:16] _7I4863_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_67 (_7I4863_$1I4488_$1I4621_SSRA, _7I4863_$1I4488_$1I4621_SSRA__vlIN);

 wire  _7I4863_$1I4488_$1I4621_SSRB;
 reg [1:16] _7I4863_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_68 (_7I4863_$1I4488_$1I4621_SSRB, _7I4863_$1I4488_$1I4621_SSRB__vlIN);

 wire  _7I4863_$1I4488_$1I4621_WEA;
 reg [1:16] _7I4863_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_69 (_7I4863_$1I4488_$1I4621_WEA, _7I4863_$1I4488_$1I4621_WEA__vlIN);

 wire  _7I4863_$1I4488_$1I4621_WEB;
 reg [1:16] _7I4863_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_70 (_7I4863_$1I4488_$1I4621_WEB, _7I4863_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _7I4863_$1I4488_$1I4621 ( _7I4863_$1I4488_$1I4621_DOA , _7I4863_$1I4488_$1I4621_DOB , _7I4863_$1I4488_$1I4621_DOPA , _7I4863_$1I4488_$1I4621_DOPB , _7I4863_$1I4488_$1I4621_ADDRA , _7I4863_$1I4488_$1I4621_ADDRB , _7I4863_$1I4488_$1I4621_CLKA , _7I4863_$1I4488_$1I4621_CLKB , _7I4863_$1I4488_$1I4621_DIA , _7I4863_$1I4488_$1I4621_DIB , _7I4863_$1I4488_$1I4621_DIPA , _7I4863_$1I4488_$1I4621_DIPB , _7I4863_$1I4488_$1I4621_ENA , _7I4863_$1I4488_$1I4621_ENB , _7I4863_$1I4488_$1I4621_SSRA , _7I4863_$1I4488_$1I4621_SSRB , _7I4863_$1I4488_$1I4621_WEA , _7I4863_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4863_$1I4488_$1I4620_DOA;

 wire [15:0] _7I4863_$1I4488_$1I4620_DOB;

 wire [0:0] _7I4863_$1I4488_$1I4620_DOPA;

 wire [1:0] _7I4863_$1I4488_$1I4620_DOPB;

 wire [10:0] _7I4863_$1I4488_$1I4620_ADDRA;
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_71_10 (_7I4863_$1I4488_$1I4620_ADDRA[10], _7I4863_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_71_9 (_7I4863_$1I4488_$1I4620_ADDRA[9], _7I4863_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_71_8 (_7I4863_$1I4488_$1I4620_ADDRA[8], _7I4863_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_71_7 (_7I4863_$1I4488_$1I4620_ADDRA[7], _7I4863_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_71_6 (_7I4863_$1I4488_$1I4620_ADDRA[6], _7I4863_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_71_5 (_7I4863_$1I4488_$1I4620_ADDRA[5], _7I4863_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_71_4 (_7I4863_$1I4488_$1I4620_ADDRA[4], _7I4863_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_71_3 (_7I4863_$1I4488_$1I4620_ADDRA[3], _7I4863_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_71_2 (_7I4863_$1I4488_$1I4620_ADDRA[2], _7I4863_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_71_1 (_7I4863_$1I4488_$1I4620_ADDRA[1], _7I4863_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_71_0 (_7I4863_$1I4488_$1I4620_ADDRA[0], _7I4863_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _7I4863_$1I4488_$1I4620_ADDRB;
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_72_9 (_7I4863_$1I4488_$1I4620_ADDRB[9], _7I4863_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_72_8 (_7I4863_$1I4488_$1I4620_ADDRB[8], _7I4863_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_72_7 (_7I4863_$1I4488_$1I4620_ADDRB[7], _7I4863_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_72_6 (_7I4863_$1I4488_$1I4620_ADDRB[6], _7I4863_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_72_5 (_7I4863_$1I4488_$1I4620_ADDRB[5], _7I4863_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_72_4 (_7I4863_$1I4488_$1I4620_ADDRB[4], _7I4863_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_72_3 (_7I4863_$1I4488_$1I4620_ADDRB[3], _7I4863_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_72_2 (_7I4863_$1I4488_$1I4620_ADDRB[2], _7I4863_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_72_1 (_7I4863_$1I4488_$1I4620_ADDRB[1], _7I4863_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_72_0 (_7I4863_$1I4488_$1I4620_ADDRB[0], _7I4863_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _7I4863_$1I4488_$1I4620_CLKA;
 reg [1:16] _7I4863_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_73 (_7I4863_$1I4488_$1I4620_CLKA, _7I4863_$1I4488_$1I4620_CLKA__vlIN);

 wire  _7I4863_$1I4488_$1I4620_CLKB;
 reg [1:16] _7I4863_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_74 (_7I4863_$1I4488_$1I4620_CLKB, _7I4863_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _7I4863_$1I4488_$1I4620_DIA;
 reg [1:16] _7I4863_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_75_7 (_7I4863_$1I4488_$1I4620_DIA[7], _7I4863_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_75_6 (_7I4863_$1I4488_$1I4620_DIA[6], _7I4863_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_75_5 (_7I4863_$1I4488_$1I4620_DIA[5], _7I4863_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_75_4 (_7I4863_$1I4488_$1I4620_DIA[4], _7I4863_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_75_3 (_7I4863_$1I4488_$1I4620_DIA[3], _7I4863_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_75_2 (_7I4863_$1I4488_$1I4620_DIA[2], _7I4863_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_75_1 (_7I4863_$1I4488_$1I4620_DIA[1], _7I4863_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_75_0 (_7I4863_$1I4488_$1I4620_DIA[0], _7I4863_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _7I4863_$1I4488_$1I4620_DIB;
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_76_15 (_7I4863_$1I4488_$1I4620_DIB[15], _7I4863_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_76_14 (_7I4863_$1I4488_$1I4620_DIB[14], _7I4863_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_76_13 (_7I4863_$1I4488_$1I4620_DIB[13], _7I4863_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_76_12 (_7I4863_$1I4488_$1I4620_DIB[12], _7I4863_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_76_11 (_7I4863_$1I4488_$1I4620_DIB[11], _7I4863_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_76_10 (_7I4863_$1I4488_$1I4620_DIB[10], _7I4863_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_76_9 (_7I4863_$1I4488_$1I4620_DIB[9], _7I4863_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_76_8 (_7I4863_$1I4488_$1I4620_DIB[8], _7I4863_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_76_7 (_7I4863_$1I4488_$1I4620_DIB[7], _7I4863_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_76_6 (_7I4863_$1I4488_$1I4620_DIB[6], _7I4863_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_76_5 (_7I4863_$1I4488_$1I4620_DIB[5], _7I4863_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_76_4 (_7I4863_$1I4488_$1I4620_DIB[4], _7I4863_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_76_3 (_7I4863_$1I4488_$1I4620_DIB[3], _7I4863_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_76_2 (_7I4863_$1I4488_$1I4620_DIB[2], _7I4863_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_76_1 (_7I4863_$1I4488_$1I4620_DIB[1], _7I4863_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_76_0 (_7I4863_$1I4488_$1I4620_DIB[0], _7I4863_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _7I4863_$1I4488_$1I4620_DIPA;
 reg [1:16] _7I4863_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_77_0 (_7I4863_$1I4488_$1I4620_DIPA[0], _7I4863_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _7I4863_$1I4488_$1I4620_DIPB;
 reg [1:16] _7I4863_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_78_1 (_7I4863_$1I4488_$1I4620_DIPB[1], _7I4863_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _7I4863_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_78_0 (_7I4863_$1I4488_$1I4620_DIPB[0], _7I4863_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _7I4863_$1I4488_$1I4620_ENA;
 reg [1:16] _7I4863_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_79 (_7I4863_$1I4488_$1I4620_ENA, _7I4863_$1I4488_$1I4620_ENA__vlIN);

 wire  _7I4863_$1I4488_$1I4620_ENB;
 reg [1:16] _7I4863_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_80 (_7I4863_$1I4488_$1I4620_ENB, _7I4863_$1I4488_$1I4620_ENB__vlIN);

 wire  _7I4863_$1I4488_$1I4620_SSRA;
 reg [1:16] _7I4863_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_81 (_7I4863_$1I4488_$1I4620_SSRA, _7I4863_$1I4488_$1I4620_SSRA__vlIN);

 wire  _7I4863_$1I4488_$1I4620_SSRB;
 reg [1:16] _7I4863_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_82 (_7I4863_$1I4488_$1I4620_SSRB, _7I4863_$1I4488_$1I4620_SSRB__vlIN);

 wire  _7I4863_$1I4488_$1I4620_WEA;
 reg [1:16] _7I4863_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_83 (_7I4863_$1I4488_$1I4620_WEA, _7I4863_$1I4488_$1I4620_WEA__vlIN);

 wire  _7I4863_$1I4488_$1I4620_WEB;
 reg [1:16] _7I4863_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_84 (_7I4863_$1I4488_$1I4620_WEB, _7I4863_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _7I4863_$1I4488_$1I4620 ( _7I4863_$1I4488_$1I4620_DOA , _7I4863_$1I4488_$1I4620_DOB , _7I4863_$1I4488_$1I4620_DOPA , _7I4863_$1I4488_$1I4620_DOPB , _7I4863_$1I4488_$1I4620_ADDRA , _7I4863_$1I4488_$1I4620_ADDRB , _7I4863_$1I4488_$1I4620_CLKA , _7I4863_$1I4488_$1I4620_CLKB , _7I4863_$1I4488_$1I4620_DIA , _7I4863_$1I4488_$1I4620_DIB , _7I4863_$1I4488_$1I4620_DIPA , _7I4863_$1I4488_$1I4620_DIPB , _7I4863_$1I4488_$1I4620_ENA , _7I4863_$1I4488_$1I4620_ENB , _7I4863_$1I4488_$1I4620_SSRA , _7I4863_$1I4488_$1I4620_SSRB , _7I4863_$1I4488_$1I4620_WEA , _7I4863_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4838_$1I4488_$1I4621_DOA;

 wire [15:0] _7I4838_$1I4488_$1I4621_DOB;

 wire [0:0] _7I4838_$1I4488_$1I4621_DOPA;

 wire [1:0] _7I4838_$1I4488_$1I4621_DOPB;

 wire [10:0] _7I4838_$1I4488_$1I4621_ADDRA;
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_85_10 (_7I4838_$1I4488_$1I4621_ADDRA[10], _7I4838_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_85_9 (_7I4838_$1I4488_$1I4621_ADDRA[9], _7I4838_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_85_8 (_7I4838_$1I4488_$1I4621_ADDRA[8], _7I4838_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_85_7 (_7I4838_$1I4488_$1I4621_ADDRA[7], _7I4838_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_85_6 (_7I4838_$1I4488_$1I4621_ADDRA[6], _7I4838_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_85_5 (_7I4838_$1I4488_$1I4621_ADDRA[5], _7I4838_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_85_4 (_7I4838_$1I4488_$1I4621_ADDRA[4], _7I4838_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_85_3 (_7I4838_$1I4488_$1I4621_ADDRA[3], _7I4838_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_85_2 (_7I4838_$1I4488_$1I4621_ADDRA[2], _7I4838_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_85_1 (_7I4838_$1I4488_$1I4621_ADDRA[1], _7I4838_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_85_0 (_7I4838_$1I4488_$1I4621_ADDRA[0], _7I4838_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _7I4838_$1I4488_$1I4621_ADDRB;
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_86_9 (_7I4838_$1I4488_$1I4621_ADDRB[9], _7I4838_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_86_8 (_7I4838_$1I4488_$1I4621_ADDRB[8], _7I4838_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_86_7 (_7I4838_$1I4488_$1I4621_ADDRB[7], _7I4838_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_86_6 (_7I4838_$1I4488_$1I4621_ADDRB[6], _7I4838_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_86_5 (_7I4838_$1I4488_$1I4621_ADDRB[5], _7I4838_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_86_4 (_7I4838_$1I4488_$1I4621_ADDRB[4], _7I4838_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_86_3 (_7I4838_$1I4488_$1I4621_ADDRB[3], _7I4838_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_86_2 (_7I4838_$1I4488_$1I4621_ADDRB[2], _7I4838_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_86_1 (_7I4838_$1I4488_$1I4621_ADDRB[1], _7I4838_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_86_0 (_7I4838_$1I4488_$1I4621_ADDRB[0], _7I4838_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _7I4838_$1I4488_$1I4621_CLKA;
 reg [1:16] _7I4838_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_87 (_7I4838_$1I4488_$1I4621_CLKA, _7I4838_$1I4488_$1I4621_CLKA__vlIN);

 wire  _7I4838_$1I4488_$1I4621_CLKB;
 reg [1:16] _7I4838_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_88 (_7I4838_$1I4488_$1I4621_CLKB, _7I4838_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _7I4838_$1I4488_$1I4621_DIA;
 reg [1:16] _7I4838_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_89_7 (_7I4838_$1I4488_$1I4621_DIA[7], _7I4838_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_89_6 (_7I4838_$1I4488_$1I4621_DIA[6], _7I4838_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_89_5 (_7I4838_$1I4488_$1I4621_DIA[5], _7I4838_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_89_4 (_7I4838_$1I4488_$1I4621_DIA[4], _7I4838_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_89_3 (_7I4838_$1I4488_$1I4621_DIA[3], _7I4838_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_89_2 (_7I4838_$1I4488_$1I4621_DIA[2], _7I4838_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_89_1 (_7I4838_$1I4488_$1I4621_DIA[1], _7I4838_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_89_0 (_7I4838_$1I4488_$1I4621_DIA[0], _7I4838_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _7I4838_$1I4488_$1I4621_DIB;
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_90_15 (_7I4838_$1I4488_$1I4621_DIB[15], _7I4838_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_90_14 (_7I4838_$1I4488_$1I4621_DIB[14], _7I4838_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_90_13 (_7I4838_$1I4488_$1I4621_DIB[13], _7I4838_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_90_12 (_7I4838_$1I4488_$1I4621_DIB[12], _7I4838_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_90_11 (_7I4838_$1I4488_$1I4621_DIB[11], _7I4838_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_90_10 (_7I4838_$1I4488_$1I4621_DIB[10], _7I4838_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_90_9 (_7I4838_$1I4488_$1I4621_DIB[9], _7I4838_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_90_8 (_7I4838_$1I4488_$1I4621_DIB[8], _7I4838_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_90_7 (_7I4838_$1I4488_$1I4621_DIB[7], _7I4838_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_90_6 (_7I4838_$1I4488_$1I4621_DIB[6], _7I4838_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_90_5 (_7I4838_$1I4488_$1I4621_DIB[5], _7I4838_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_90_4 (_7I4838_$1I4488_$1I4621_DIB[4], _7I4838_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_90_3 (_7I4838_$1I4488_$1I4621_DIB[3], _7I4838_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_90_2 (_7I4838_$1I4488_$1I4621_DIB[2], _7I4838_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_90_1 (_7I4838_$1I4488_$1I4621_DIB[1], _7I4838_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_90_0 (_7I4838_$1I4488_$1I4621_DIB[0], _7I4838_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _7I4838_$1I4488_$1I4621_DIPA;
 reg [1:16] _7I4838_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_91_0 (_7I4838_$1I4488_$1I4621_DIPA[0], _7I4838_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _7I4838_$1I4488_$1I4621_DIPB;
 reg [1:16] _7I4838_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_92_1 (_7I4838_$1I4488_$1I4621_DIPB[1], _7I4838_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_92_0 (_7I4838_$1I4488_$1I4621_DIPB[0], _7I4838_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _7I4838_$1I4488_$1I4621_ENA;
 reg [1:16] _7I4838_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_93 (_7I4838_$1I4488_$1I4621_ENA, _7I4838_$1I4488_$1I4621_ENA__vlIN);

 wire  _7I4838_$1I4488_$1I4621_ENB;
 reg [1:16] _7I4838_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_94 (_7I4838_$1I4488_$1I4621_ENB, _7I4838_$1I4488_$1I4621_ENB__vlIN);

 wire  _7I4838_$1I4488_$1I4621_SSRA;
 reg [1:16] _7I4838_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_95 (_7I4838_$1I4488_$1I4621_SSRA, _7I4838_$1I4488_$1I4621_SSRA__vlIN);

 wire  _7I4838_$1I4488_$1I4621_SSRB;
 reg [1:16] _7I4838_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_96 (_7I4838_$1I4488_$1I4621_SSRB, _7I4838_$1I4488_$1I4621_SSRB__vlIN);

 wire  _7I4838_$1I4488_$1I4621_WEA;
 reg [1:16] _7I4838_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_97 (_7I4838_$1I4488_$1I4621_WEA, _7I4838_$1I4488_$1I4621_WEA__vlIN);

 wire  _7I4838_$1I4488_$1I4621_WEB;
 reg [1:16] _7I4838_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_98 (_7I4838_$1I4488_$1I4621_WEB, _7I4838_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _7I4838_$1I4488_$1I4621 ( _7I4838_$1I4488_$1I4621_DOA , _7I4838_$1I4488_$1I4621_DOB , _7I4838_$1I4488_$1I4621_DOPA , _7I4838_$1I4488_$1I4621_DOPB , _7I4838_$1I4488_$1I4621_ADDRA , _7I4838_$1I4488_$1I4621_ADDRB , _7I4838_$1I4488_$1I4621_CLKA , _7I4838_$1I4488_$1I4621_CLKB , _7I4838_$1I4488_$1I4621_DIA , _7I4838_$1I4488_$1I4621_DIB , _7I4838_$1I4488_$1I4621_DIPA , _7I4838_$1I4488_$1I4621_DIPB , _7I4838_$1I4488_$1I4621_ENA , _7I4838_$1I4488_$1I4621_ENB , _7I4838_$1I4488_$1I4621_SSRA , _7I4838_$1I4488_$1I4621_SSRB , _7I4838_$1I4488_$1I4621_WEA , _7I4838_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4838_$1I4488_$1I4620_DOA;

 wire [15:0] _7I4838_$1I4488_$1I4620_DOB;

 wire [0:0] _7I4838_$1I4488_$1I4620_DOPA;

 wire [1:0] _7I4838_$1I4488_$1I4620_DOPB;

 wire [10:0] _7I4838_$1I4488_$1I4620_ADDRA;
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_99_10 (_7I4838_$1I4488_$1I4620_ADDRA[10], _7I4838_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_99_9 (_7I4838_$1I4488_$1I4620_ADDRA[9], _7I4838_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_99_8 (_7I4838_$1I4488_$1I4620_ADDRA[8], _7I4838_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_99_7 (_7I4838_$1I4488_$1I4620_ADDRA[7], _7I4838_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_99_6 (_7I4838_$1I4488_$1I4620_ADDRA[6], _7I4838_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_99_5 (_7I4838_$1I4488_$1I4620_ADDRA[5], _7I4838_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_99_4 (_7I4838_$1I4488_$1I4620_ADDRA[4], _7I4838_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_99_3 (_7I4838_$1I4488_$1I4620_ADDRA[3], _7I4838_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_99_2 (_7I4838_$1I4488_$1I4620_ADDRA[2], _7I4838_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_99_1 (_7I4838_$1I4488_$1I4620_ADDRA[1], _7I4838_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_99_0 (_7I4838_$1I4488_$1I4620_ADDRA[0], _7I4838_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _7I4838_$1I4488_$1I4620_ADDRB;
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_100_9 (_7I4838_$1I4488_$1I4620_ADDRB[9], _7I4838_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_100_8 (_7I4838_$1I4488_$1I4620_ADDRB[8], _7I4838_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_100_7 (_7I4838_$1I4488_$1I4620_ADDRB[7], _7I4838_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_100_6 (_7I4838_$1I4488_$1I4620_ADDRB[6], _7I4838_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_100_5 (_7I4838_$1I4488_$1I4620_ADDRB[5], _7I4838_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_100_4 (_7I4838_$1I4488_$1I4620_ADDRB[4], _7I4838_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_100_3 (_7I4838_$1I4488_$1I4620_ADDRB[3], _7I4838_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_100_2 (_7I4838_$1I4488_$1I4620_ADDRB[2], _7I4838_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_100_1 (_7I4838_$1I4488_$1I4620_ADDRB[1], _7I4838_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_100_0 (_7I4838_$1I4488_$1I4620_ADDRB[0], _7I4838_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _7I4838_$1I4488_$1I4620_CLKA;
 reg [1:16] _7I4838_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_101 (_7I4838_$1I4488_$1I4620_CLKA, _7I4838_$1I4488_$1I4620_CLKA__vlIN);

 wire  _7I4838_$1I4488_$1I4620_CLKB;
 reg [1:16] _7I4838_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_102 (_7I4838_$1I4488_$1I4620_CLKB, _7I4838_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _7I4838_$1I4488_$1I4620_DIA;
 reg [1:16] _7I4838_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_103_7 (_7I4838_$1I4488_$1I4620_DIA[7], _7I4838_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_103_6 (_7I4838_$1I4488_$1I4620_DIA[6], _7I4838_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_103_5 (_7I4838_$1I4488_$1I4620_DIA[5], _7I4838_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_103_4 (_7I4838_$1I4488_$1I4620_DIA[4], _7I4838_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_103_3 (_7I4838_$1I4488_$1I4620_DIA[3], _7I4838_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_103_2 (_7I4838_$1I4488_$1I4620_DIA[2], _7I4838_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_103_1 (_7I4838_$1I4488_$1I4620_DIA[1], _7I4838_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_103_0 (_7I4838_$1I4488_$1I4620_DIA[0], _7I4838_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _7I4838_$1I4488_$1I4620_DIB;
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_104_15 (_7I4838_$1I4488_$1I4620_DIB[15], _7I4838_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_104_14 (_7I4838_$1I4488_$1I4620_DIB[14], _7I4838_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_104_13 (_7I4838_$1I4488_$1I4620_DIB[13], _7I4838_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_104_12 (_7I4838_$1I4488_$1I4620_DIB[12], _7I4838_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_104_11 (_7I4838_$1I4488_$1I4620_DIB[11], _7I4838_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_104_10 (_7I4838_$1I4488_$1I4620_DIB[10], _7I4838_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_104_9 (_7I4838_$1I4488_$1I4620_DIB[9], _7I4838_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_104_8 (_7I4838_$1I4488_$1I4620_DIB[8], _7I4838_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_104_7 (_7I4838_$1I4488_$1I4620_DIB[7], _7I4838_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_104_6 (_7I4838_$1I4488_$1I4620_DIB[6], _7I4838_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_104_5 (_7I4838_$1I4488_$1I4620_DIB[5], _7I4838_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_104_4 (_7I4838_$1I4488_$1I4620_DIB[4], _7I4838_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_104_3 (_7I4838_$1I4488_$1I4620_DIB[3], _7I4838_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_104_2 (_7I4838_$1I4488_$1I4620_DIB[2], _7I4838_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_104_1 (_7I4838_$1I4488_$1I4620_DIB[1], _7I4838_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_104_0 (_7I4838_$1I4488_$1I4620_DIB[0], _7I4838_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _7I4838_$1I4488_$1I4620_DIPA;
 reg [1:16] _7I4838_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_105_0 (_7I4838_$1I4488_$1I4620_DIPA[0], _7I4838_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _7I4838_$1I4488_$1I4620_DIPB;
 reg [1:16] _7I4838_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_106_1 (_7I4838_$1I4488_$1I4620_DIPB[1], _7I4838_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _7I4838_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_106_0 (_7I4838_$1I4488_$1I4620_DIPB[0], _7I4838_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _7I4838_$1I4488_$1I4620_ENA;
 reg [1:16] _7I4838_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_107 (_7I4838_$1I4488_$1I4620_ENA, _7I4838_$1I4488_$1I4620_ENA__vlIN);

 wire  _7I4838_$1I4488_$1I4620_ENB;
 reg [1:16] _7I4838_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_108 (_7I4838_$1I4488_$1I4620_ENB, _7I4838_$1I4488_$1I4620_ENB__vlIN);

 wire  _7I4838_$1I4488_$1I4620_SSRA;
 reg [1:16] _7I4838_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_109 (_7I4838_$1I4488_$1I4620_SSRA, _7I4838_$1I4488_$1I4620_SSRA__vlIN);

 wire  _7I4838_$1I4488_$1I4620_SSRB;
 reg [1:16] _7I4838_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_110 (_7I4838_$1I4488_$1I4620_SSRB, _7I4838_$1I4488_$1I4620_SSRB__vlIN);

 wire  _7I4838_$1I4488_$1I4620_WEA;
 reg [1:16] _7I4838_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_111 (_7I4838_$1I4488_$1I4620_WEA, _7I4838_$1I4488_$1I4620_WEA__vlIN);

 wire  _7I4838_$1I4488_$1I4620_WEB;
 reg [1:16] _7I4838_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_112 (_7I4838_$1I4488_$1I4620_WEB, _7I4838_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _7I4838_$1I4488_$1I4620 ( _7I4838_$1I4488_$1I4620_DOA , _7I4838_$1I4488_$1I4620_DOB , _7I4838_$1I4488_$1I4620_DOPA , _7I4838_$1I4488_$1I4620_DOPB , _7I4838_$1I4488_$1I4620_ADDRA , _7I4838_$1I4488_$1I4620_ADDRB , _7I4838_$1I4488_$1I4620_CLKA , _7I4838_$1I4488_$1I4620_CLKB , _7I4838_$1I4488_$1I4620_DIA , _7I4838_$1I4488_$1I4620_DIB , _7I4838_$1I4488_$1I4620_DIPA , _7I4838_$1I4488_$1I4620_DIPB , _7I4838_$1I4488_$1I4620_ENA , _7I4838_$1I4488_$1I4620_ENB , _7I4838_$1I4488_$1I4620_SSRA , _7I4838_$1I4488_$1I4620_SSRB , _7I4838_$1I4488_$1I4620_WEA , _7I4838_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4762_$1I4488_$1I4621_DOA;

 wire [15:0] _7I4762_$1I4488_$1I4621_DOB;

 wire [0:0] _7I4762_$1I4488_$1I4621_DOPA;

 wire [1:0] _7I4762_$1I4488_$1I4621_DOPB;

 wire [10:0] _7I4762_$1I4488_$1I4621_ADDRA;
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_113_10 (_7I4762_$1I4488_$1I4621_ADDRA[10], _7I4762_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_113_9 (_7I4762_$1I4488_$1I4621_ADDRA[9], _7I4762_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_113_8 (_7I4762_$1I4488_$1I4621_ADDRA[8], _7I4762_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_113_7 (_7I4762_$1I4488_$1I4621_ADDRA[7], _7I4762_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_113_6 (_7I4762_$1I4488_$1I4621_ADDRA[6], _7I4762_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_113_5 (_7I4762_$1I4488_$1I4621_ADDRA[5], _7I4762_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_113_4 (_7I4762_$1I4488_$1I4621_ADDRA[4], _7I4762_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_113_3 (_7I4762_$1I4488_$1I4621_ADDRA[3], _7I4762_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_113_2 (_7I4762_$1I4488_$1I4621_ADDRA[2], _7I4762_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_113_1 (_7I4762_$1I4488_$1I4621_ADDRA[1], _7I4762_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_113_0 (_7I4762_$1I4488_$1I4621_ADDRA[0], _7I4762_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _7I4762_$1I4488_$1I4621_ADDRB;
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_114_9 (_7I4762_$1I4488_$1I4621_ADDRB[9], _7I4762_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_114_8 (_7I4762_$1I4488_$1I4621_ADDRB[8], _7I4762_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_114_7 (_7I4762_$1I4488_$1I4621_ADDRB[7], _7I4762_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_114_6 (_7I4762_$1I4488_$1I4621_ADDRB[6], _7I4762_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_114_5 (_7I4762_$1I4488_$1I4621_ADDRB[5], _7I4762_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_114_4 (_7I4762_$1I4488_$1I4621_ADDRB[4], _7I4762_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_114_3 (_7I4762_$1I4488_$1I4621_ADDRB[3], _7I4762_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_114_2 (_7I4762_$1I4488_$1I4621_ADDRB[2], _7I4762_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_114_1 (_7I4762_$1I4488_$1I4621_ADDRB[1], _7I4762_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_114_0 (_7I4762_$1I4488_$1I4621_ADDRB[0], _7I4762_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _7I4762_$1I4488_$1I4621_CLKA;
 reg [1:16] _7I4762_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_115 (_7I4762_$1I4488_$1I4621_CLKA, _7I4762_$1I4488_$1I4621_CLKA__vlIN);

 wire  _7I4762_$1I4488_$1I4621_CLKB;
 reg [1:16] _7I4762_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_116 (_7I4762_$1I4488_$1I4621_CLKB, _7I4762_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _7I4762_$1I4488_$1I4621_DIA;
 reg [1:16] _7I4762_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_117_7 (_7I4762_$1I4488_$1I4621_DIA[7], _7I4762_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_117_6 (_7I4762_$1I4488_$1I4621_DIA[6], _7I4762_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_117_5 (_7I4762_$1I4488_$1I4621_DIA[5], _7I4762_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_117_4 (_7I4762_$1I4488_$1I4621_DIA[4], _7I4762_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_117_3 (_7I4762_$1I4488_$1I4621_DIA[3], _7I4762_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_117_2 (_7I4762_$1I4488_$1I4621_DIA[2], _7I4762_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_117_1 (_7I4762_$1I4488_$1I4621_DIA[1], _7I4762_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_117_0 (_7I4762_$1I4488_$1I4621_DIA[0], _7I4762_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _7I4762_$1I4488_$1I4621_DIB;
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_118_15 (_7I4762_$1I4488_$1I4621_DIB[15], _7I4762_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_118_14 (_7I4762_$1I4488_$1I4621_DIB[14], _7I4762_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_118_13 (_7I4762_$1I4488_$1I4621_DIB[13], _7I4762_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_118_12 (_7I4762_$1I4488_$1I4621_DIB[12], _7I4762_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_118_11 (_7I4762_$1I4488_$1I4621_DIB[11], _7I4762_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_118_10 (_7I4762_$1I4488_$1I4621_DIB[10], _7I4762_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_118_9 (_7I4762_$1I4488_$1I4621_DIB[9], _7I4762_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_118_8 (_7I4762_$1I4488_$1I4621_DIB[8], _7I4762_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_118_7 (_7I4762_$1I4488_$1I4621_DIB[7], _7I4762_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_118_6 (_7I4762_$1I4488_$1I4621_DIB[6], _7I4762_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_118_5 (_7I4762_$1I4488_$1I4621_DIB[5], _7I4762_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_118_4 (_7I4762_$1I4488_$1I4621_DIB[4], _7I4762_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_118_3 (_7I4762_$1I4488_$1I4621_DIB[3], _7I4762_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_118_2 (_7I4762_$1I4488_$1I4621_DIB[2], _7I4762_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_118_1 (_7I4762_$1I4488_$1I4621_DIB[1], _7I4762_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_118_0 (_7I4762_$1I4488_$1I4621_DIB[0], _7I4762_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _7I4762_$1I4488_$1I4621_DIPA;
 reg [1:16] _7I4762_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_119_0 (_7I4762_$1I4488_$1I4621_DIPA[0], _7I4762_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _7I4762_$1I4488_$1I4621_DIPB;
 reg [1:16] _7I4762_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_120_1 (_7I4762_$1I4488_$1I4621_DIPB[1], _7I4762_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_120_0 (_7I4762_$1I4488_$1I4621_DIPB[0], _7I4762_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _7I4762_$1I4488_$1I4621_ENA;
 reg [1:16] _7I4762_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_121 (_7I4762_$1I4488_$1I4621_ENA, _7I4762_$1I4488_$1I4621_ENA__vlIN);

 wire  _7I4762_$1I4488_$1I4621_ENB;
 reg [1:16] _7I4762_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_122 (_7I4762_$1I4488_$1I4621_ENB, _7I4762_$1I4488_$1I4621_ENB__vlIN);

 wire  _7I4762_$1I4488_$1I4621_SSRA;
 reg [1:16] _7I4762_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_123 (_7I4762_$1I4488_$1I4621_SSRA, _7I4762_$1I4488_$1I4621_SSRA__vlIN);

 wire  _7I4762_$1I4488_$1I4621_SSRB;
 reg [1:16] _7I4762_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_124 (_7I4762_$1I4488_$1I4621_SSRB, _7I4762_$1I4488_$1I4621_SSRB__vlIN);

 wire  _7I4762_$1I4488_$1I4621_WEA;
 reg [1:16] _7I4762_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_125 (_7I4762_$1I4488_$1I4621_WEA, _7I4762_$1I4488_$1I4621_WEA__vlIN);

 wire  _7I4762_$1I4488_$1I4621_WEB;
 reg [1:16] _7I4762_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_126 (_7I4762_$1I4488_$1I4621_WEB, _7I4762_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _7I4762_$1I4488_$1I4621 ( _7I4762_$1I4488_$1I4621_DOA , _7I4762_$1I4488_$1I4621_DOB , _7I4762_$1I4488_$1I4621_DOPA , _7I4762_$1I4488_$1I4621_DOPB , _7I4762_$1I4488_$1I4621_ADDRA , _7I4762_$1I4488_$1I4621_ADDRB , _7I4762_$1I4488_$1I4621_CLKA , _7I4762_$1I4488_$1I4621_CLKB , _7I4762_$1I4488_$1I4621_DIA , _7I4762_$1I4488_$1I4621_DIB , _7I4762_$1I4488_$1I4621_DIPA , _7I4762_$1I4488_$1I4621_DIPB , _7I4762_$1I4488_$1I4621_ENA , _7I4762_$1I4488_$1I4621_ENB , _7I4762_$1I4488_$1I4621_SSRA , _7I4762_$1I4488_$1I4621_SSRB , _7I4762_$1I4488_$1I4621_WEA , _7I4762_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4762_$1I4488_$1I4620_DOA;

 wire [15:0] _7I4762_$1I4488_$1I4620_DOB;

 wire [0:0] _7I4762_$1I4488_$1I4620_DOPA;

 wire [1:0] _7I4762_$1I4488_$1I4620_DOPB;

 wire [10:0] _7I4762_$1I4488_$1I4620_ADDRA;
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_127_10 (_7I4762_$1I4488_$1I4620_ADDRA[10], _7I4762_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_127_9 (_7I4762_$1I4488_$1I4620_ADDRA[9], _7I4762_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_127_8 (_7I4762_$1I4488_$1I4620_ADDRA[8], _7I4762_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_127_7 (_7I4762_$1I4488_$1I4620_ADDRA[7], _7I4762_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_127_6 (_7I4762_$1I4488_$1I4620_ADDRA[6], _7I4762_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_127_5 (_7I4762_$1I4488_$1I4620_ADDRA[5], _7I4762_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_127_4 (_7I4762_$1I4488_$1I4620_ADDRA[4], _7I4762_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_127_3 (_7I4762_$1I4488_$1I4620_ADDRA[3], _7I4762_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_127_2 (_7I4762_$1I4488_$1I4620_ADDRA[2], _7I4762_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_127_1 (_7I4762_$1I4488_$1I4620_ADDRA[1], _7I4762_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_127_0 (_7I4762_$1I4488_$1I4620_ADDRA[0], _7I4762_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _7I4762_$1I4488_$1I4620_ADDRB;
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_128_9 (_7I4762_$1I4488_$1I4620_ADDRB[9], _7I4762_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_128_8 (_7I4762_$1I4488_$1I4620_ADDRB[8], _7I4762_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_128_7 (_7I4762_$1I4488_$1I4620_ADDRB[7], _7I4762_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_128_6 (_7I4762_$1I4488_$1I4620_ADDRB[6], _7I4762_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_128_5 (_7I4762_$1I4488_$1I4620_ADDRB[5], _7I4762_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_128_4 (_7I4762_$1I4488_$1I4620_ADDRB[4], _7I4762_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_128_3 (_7I4762_$1I4488_$1I4620_ADDRB[3], _7I4762_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_128_2 (_7I4762_$1I4488_$1I4620_ADDRB[2], _7I4762_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_128_1 (_7I4762_$1I4488_$1I4620_ADDRB[1], _7I4762_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_128_0 (_7I4762_$1I4488_$1I4620_ADDRB[0], _7I4762_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _7I4762_$1I4488_$1I4620_CLKA;
 reg [1:16] _7I4762_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_129 (_7I4762_$1I4488_$1I4620_CLKA, _7I4762_$1I4488_$1I4620_CLKA__vlIN);

 wire  _7I4762_$1I4488_$1I4620_CLKB;
 reg [1:16] _7I4762_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_130 (_7I4762_$1I4488_$1I4620_CLKB, _7I4762_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _7I4762_$1I4488_$1I4620_DIA;
 reg [1:16] _7I4762_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_131_7 (_7I4762_$1I4488_$1I4620_DIA[7], _7I4762_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_131_6 (_7I4762_$1I4488_$1I4620_DIA[6], _7I4762_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_131_5 (_7I4762_$1I4488_$1I4620_DIA[5], _7I4762_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_131_4 (_7I4762_$1I4488_$1I4620_DIA[4], _7I4762_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_131_3 (_7I4762_$1I4488_$1I4620_DIA[3], _7I4762_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_131_2 (_7I4762_$1I4488_$1I4620_DIA[2], _7I4762_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_131_1 (_7I4762_$1I4488_$1I4620_DIA[1], _7I4762_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_131_0 (_7I4762_$1I4488_$1I4620_DIA[0], _7I4762_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _7I4762_$1I4488_$1I4620_DIB;
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_132_15 (_7I4762_$1I4488_$1I4620_DIB[15], _7I4762_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_132_14 (_7I4762_$1I4488_$1I4620_DIB[14], _7I4762_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_132_13 (_7I4762_$1I4488_$1I4620_DIB[13], _7I4762_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_132_12 (_7I4762_$1I4488_$1I4620_DIB[12], _7I4762_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_132_11 (_7I4762_$1I4488_$1I4620_DIB[11], _7I4762_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_132_10 (_7I4762_$1I4488_$1I4620_DIB[10], _7I4762_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_132_9 (_7I4762_$1I4488_$1I4620_DIB[9], _7I4762_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_132_8 (_7I4762_$1I4488_$1I4620_DIB[8], _7I4762_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_132_7 (_7I4762_$1I4488_$1I4620_DIB[7], _7I4762_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_132_6 (_7I4762_$1I4488_$1I4620_DIB[6], _7I4762_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_132_5 (_7I4762_$1I4488_$1I4620_DIB[5], _7I4762_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_132_4 (_7I4762_$1I4488_$1I4620_DIB[4], _7I4762_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_132_3 (_7I4762_$1I4488_$1I4620_DIB[3], _7I4762_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_132_2 (_7I4762_$1I4488_$1I4620_DIB[2], _7I4762_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_132_1 (_7I4762_$1I4488_$1I4620_DIB[1], _7I4762_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_132_0 (_7I4762_$1I4488_$1I4620_DIB[0], _7I4762_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _7I4762_$1I4488_$1I4620_DIPA;
 reg [1:16] _7I4762_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_133_0 (_7I4762_$1I4488_$1I4620_DIPA[0], _7I4762_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _7I4762_$1I4488_$1I4620_DIPB;
 reg [1:16] _7I4762_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_134_1 (_7I4762_$1I4488_$1I4620_DIPB[1], _7I4762_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _7I4762_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_134_0 (_7I4762_$1I4488_$1I4620_DIPB[0], _7I4762_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _7I4762_$1I4488_$1I4620_ENA;
 reg [1:16] _7I4762_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_135 (_7I4762_$1I4488_$1I4620_ENA, _7I4762_$1I4488_$1I4620_ENA__vlIN);

 wire  _7I4762_$1I4488_$1I4620_ENB;
 reg [1:16] _7I4762_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_136 (_7I4762_$1I4488_$1I4620_ENB, _7I4762_$1I4488_$1I4620_ENB__vlIN);

 wire  _7I4762_$1I4488_$1I4620_SSRA;
 reg [1:16] _7I4762_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_137 (_7I4762_$1I4488_$1I4620_SSRA, _7I4762_$1I4488_$1I4620_SSRA__vlIN);

 wire  _7I4762_$1I4488_$1I4620_SSRB;
 reg [1:16] _7I4762_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_138 (_7I4762_$1I4488_$1I4620_SSRB, _7I4762_$1I4488_$1I4620_SSRB__vlIN);

 wire  _7I4762_$1I4488_$1I4620_WEA;
 reg [1:16] _7I4762_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_139 (_7I4762_$1I4488_$1I4620_WEA, _7I4762_$1I4488_$1I4620_WEA__vlIN);

 wire  _7I4762_$1I4488_$1I4620_WEB;
 reg [1:16] _7I4762_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_140 (_7I4762_$1I4488_$1I4620_WEB, _7I4762_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _7I4762_$1I4488_$1I4620 ( _7I4762_$1I4488_$1I4620_DOA , _7I4762_$1I4488_$1I4620_DOB , _7I4762_$1I4488_$1I4620_DOPA , _7I4762_$1I4488_$1I4620_DOPB , _7I4762_$1I4488_$1I4620_ADDRA , _7I4762_$1I4488_$1I4620_ADDRB , _7I4762_$1I4488_$1I4620_CLKA , _7I4762_$1I4488_$1I4620_CLKB , _7I4762_$1I4488_$1I4620_DIA , _7I4762_$1I4488_$1I4620_DIB , _7I4762_$1I4488_$1I4620_DIPA , _7I4762_$1I4488_$1I4620_DIPB , _7I4762_$1I4488_$1I4620_ENA , _7I4762_$1I4488_$1I4620_ENB , _7I4762_$1I4488_$1I4620_SSRA , _7I4762_$1I4488_$1I4620_SSRB , _7I4762_$1I4488_$1I4620_WEA , _7I4762_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4731_$1I4488_$1I4621_DOA;

 wire [15:0] _7I4731_$1I4488_$1I4621_DOB;

 wire [0:0] _7I4731_$1I4488_$1I4621_DOPA;

 wire [1:0] _7I4731_$1I4488_$1I4621_DOPB;

 wire [10:0] _7I4731_$1I4488_$1I4621_ADDRA;
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_141_10 (_7I4731_$1I4488_$1I4621_ADDRA[10], _7I4731_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_141_9 (_7I4731_$1I4488_$1I4621_ADDRA[9], _7I4731_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_141_8 (_7I4731_$1I4488_$1I4621_ADDRA[8], _7I4731_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_141_7 (_7I4731_$1I4488_$1I4621_ADDRA[7], _7I4731_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_141_6 (_7I4731_$1I4488_$1I4621_ADDRA[6], _7I4731_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_141_5 (_7I4731_$1I4488_$1I4621_ADDRA[5], _7I4731_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_141_4 (_7I4731_$1I4488_$1I4621_ADDRA[4], _7I4731_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_141_3 (_7I4731_$1I4488_$1I4621_ADDRA[3], _7I4731_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_141_2 (_7I4731_$1I4488_$1I4621_ADDRA[2], _7I4731_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_141_1 (_7I4731_$1I4488_$1I4621_ADDRA[1], _7I4731_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_141_0 (_7I4731_$1I4488_$1I4621_ADDRA[0], _7I4731_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _7I4731_$1I4488_$1I4621_ADDRB;
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_142_9 (_7I4731_$1I4488_$1I4621_ADDRB[9], _7I4731_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_142_8 (_7I4731_$1I4488_$1I4621_ADDRB[8], _7I4731_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_142_7 (_7I4731_$1I4488_$1I4621_ADDRB[7], _7I4731_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_142_6 (_7I4731_$1I4488_$1I4621_ADDRB[6], _7I4731_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_142_5 (_7I4731_$1I4488_$1I4621_ADDRB[5], _7I4731_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_142_4 (_7I4731_$1I4488_$1I4621_ADDRB[4], _7I4731_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_142_3 (_7I4731_$1I4488_$1I4621_ADDRB[3], _7I4731_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_142_2 (_7I4731_$1I4488_$1I4621_ADDRB[2], _7I4731_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_142_1 (_7I4731_$1I4488_$1I4621_ADDRB[1], _7I4731_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_142_0 (_7I4731_$1I4488_$1I4621_ADDRB[0], _7I4731_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _7I4731_$1I4488_$1I4621_CLKA;
 reg [1:16] _7I4731_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_143 (_7I4731_$1I4488_$1I4621_CLKA, _7I4731_$1I4488_$1I4621_CLKA__vlIN);

 wire  _7I4731_$1I4488_$1I4621_CLKB;
 reg [1:16] _7I4731_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_144 (_7I4731_$1I4488_$1I4621_CLKB, _7I4731_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _7I4731_$1I4488_$1I4621_DIA;
 reg [1:16] _7I4731_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_145_7 (_7I4731_$1I4488_$1I4621_DIA[7], _7I4731_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_145_6 (_7I4731_$1I4488_$1I4621_DIA[6], _7I4731_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_145_5 (_7I4731_$1I4488_$1I4621_DIA[5], _7I4731_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_145_4 (_7I4731_$1I4488_$1I4621_DIA[4], _7I4731_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_145_3 (_7I4731_$1I4488_$1I4621_DIA[3], _7I4731_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_145_2 (_7I4731_$1I4488_$1I4621_DIA[2], _7I4731_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_145_1 (_7I4731_$1I4488_$1I4621_DIA[1], _7I4731_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_145_0 (_7I4731_$1I4488_$1I4621_DIA[0], _7I4731_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _7I4731_$1I4488_$1I4621_DIB;
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_146_15 (_7I4731_$1I4488_$1I4621_DIB[15], _7I4731_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_146_14 (_7I4731_$1I4488_$1I4621_DIB[14], _7I4731_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_146_13 (_7I4731_$1I4488_$1I4621_DIB[13], _7I4731_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_146_12 (_7I4731_$1I4488_$1I4621_DIB[12], _7I4731_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_146_11 (_7I4731_$1I4488_$1I4621_DIB[11], _7I4731_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_146_10 (_7I4731_$1I4488_$1I4621_DIB[10], _7I4731_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_146_9 (_7I4731_$1I4488_$1I4621_DIB[9], _7I4731_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_146_8 (_7I4731_$1I4488_$1I4621_DIB[8], _7I4731_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_146_7 (_7I4731_$1I4488_$1I4621_DIB[7], _7I4731_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_146_6 (_7I4731_$1I4488_$1I4621_DIB[6], _7I4731_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_146_5 (_7I4731_$1I4488_$1I4621_DIB[5], _7I4731_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_146_4 (_7I4731_$1I4488_$1I4621_DIB[4], _7I4731_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_146_3 (_7I4731_$1I4488_$1I4621_DIB[3], _7I4731_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_146_2 (_7I4731_$1I4488_$1I4621_DIB[2], _7I4731_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_146_1 (_7I4731_$1I4488_$1I4621_DIB[1], _7I4731_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_146_0 (_7I4731_$1I4488_$1I4621_DIB[0], _7I4731_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _7I4731_$1I4488_$1I4621_DIPA;
 reg [1:16] _7I4731_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_147_0 (_7I4731_$1I4488_$1I4621_DIPA[0], _7I4731_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _7I4731_$1I4488_$1I4621_DIPB;
 reg [1:16] _7I4731_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_148_1 (_7I4731_$1I4488_$1I4621_DIPB[1], _7I4731_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_148_0 (_7I4731_$1I4488_$1I4621_DIPB[0], _7I4731_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _7I4731_$1I4488_$1I4621_ENA;
 reg [1:16] _7I4731_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_149 (_7I4731_$1I4488_$1I4621_ENA, _7I4731_$1I4488_$1I4621_ENA__vlIN);

 wire  _7I4731_$1I4488_$1I4621_ENB;
 reg [1:16] _7I4731_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_150 (_7I4731_$1I4488_$1I4621_ENB, _7I4731_$1I4488_$1I4621_ENB__vlIN);

 wire  _7I4731_$1I4488_$1I4621_SSRA;
 reg [1:16] _7I4731_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_151 (_7I4731_$1I4488_$1I4621_SSRA, _7I4731_$1I4488_$1I4621_SSRA__vlIN);

 wire  _7I4731_$1I4488_$1I4621_SSRB;
 reg [1:16] _7I4731_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_152 (_7I4731_$1I4488_$1I4621_SSRB, _7I4731_$1I4488_$1I4621_SSRB__vlIN);

 wire  _7I4731_$1I4488_$1I4621_WEA;
 reg [1:16] _7I4731_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_153 (_7I4731_$1I4488_$1I4621_WEA, _7I4731_$1I4488_$1I4621_WEA__vlIN);

 wire  _7I4731_$1I4488_$1I4621_WEB;
 reg [1:16] _7I4731_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_154 (_7I4731_$1I4488_$1I4621_WEB, _7I4731_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _7I4731_$1I4488_$1I4621 ( _7I4731_$1I4488_$1I4621_DOA , _7I4731_$1I4488_$1I4621_DOB , _7I4731_$1I4488_$1I4621_DOPA , _7I4731_$1I4488_$1I4621_DOPB , _7I4731_$1I4488_$1I4621_ADDRA , _7I4731_$1I4488_$1I4621_ADDRB , _7I4731_$1I4488_$1I4621_CLKA , _7I4731_$1I4488_$1I4621_CLKB , _7I4731_$1I4488_$1I4621_DIA , _7I4731_$1I4488_$1I4621_DIB , _7I4731_$1I4488_$1I4621_DIPA , _7I4731_$1I4488_$1I4621_DIPB , _7I4731_$1I4488_$1I4621_ENA , _7I4731_$1I4488_$1I4621_ENB , _7I4731_$1I4488_$1I4621_SSRA , _7I4731_$1I4488_$1I4621_SSRB , _7I4731_$1I4488_$1I4621_WEA , _7I4731_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4731_$1I4488_$1I4620_DOA;

 wire [15:0] _7I4731_$1I4488_$1I4620_DOB;

 wire [0:0] _7I4731_$1I4488_$1I4620_DOPA;

 wire [1:0] _7I4731_$1I4488_$1I4620_DOPB;

 wire [10:0] _7I4731_$1I4488_$1I4620_ADDRA;
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_155_10 (_7I4731_$1I4488_$1I4620_ADDRA[10], _7I4731_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_155_9 (_7I4731_$1I4488_$1I4620_ADDRA[9], _7I4731_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_155_8 (_7I4731_$1I4488_$1I4620_ADDRA[8], _7I4731_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_155_7 (_7I4731_$1I4488_$1I4620_ADDRA[7], _7I4731_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_155_6 (_7I4731_$1I4488_$1I4620_ADDRA[6], _7I4731_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_155_5 (_7I4731_$1I4488_$1I4620_ADDRA[5], _7I4731_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_155_4 (_7I4731_$1I4488_$1I4620_ADDRA[4], _7I4731_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_155_3 (_7I4731_$1I4488_$1I4620_ADDRA[3], _7I4731_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_155_2 (_7I4731_$1I4488_$1I4620_ADDRA[2], _7I4731_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_155_1 (_7I4731_$1I4488_$1I4620_ADDRA[1], _7I4731_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_155_0 (_7I4731_$1I4488_$1I4620_ADDRA[0], _7I4731_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _7I4731_$1I4488_$1I4620_ADDRB;
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_156_9 (_7I4731_$1I4488_$1I4620_ADDRB[9], _7I4731_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_156_8 (_7I4731_$1I4488_$1I4620_ADDRB[8], _7I4731_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_156_7 (_7I4731_$1I4488_$1I4620_ADDRB[7], _7I4731_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_156_6 (_7I4731_$1I4488_$1I4620_ADDRB[6], _7I4731_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_156_5 (_7I4731_$1I4488_$1I4620_ADDRB[5], _7I4731_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_156_4 (_7I4731_$1I4488_$1I4620_ADDRB[4], _7I4731_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_156_3 (_7I4731_$1I4488_$1I4620_ADDRB[3], _7I4731_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_156_2 (_7I4731_$1I4488_$1I4620_ADDRB[2], _7I4731_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_156_1 (_7I4731_$1I4488_$1I4620_ADDRB[1], _7I4731_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_156_0 (_7I4731_$1I4488_$1I4620_ADDRB[0], _7I4731_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _7I4731_$1I4488_$1I4620_CLKA;
 reg [1:16] _7I4731_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_157 (_7I4731_$1I4488_$1I4620_CLKA, _7I4731_$1I4488_$1I4620_CLKA__vlIN);

 wire  _7I4731_$1I4488_$1I4620_CLKB;
 reg [1:16] _7I4731_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_158 (_7I4731_$1I4488_$1I4620_CLKB, _7I4731_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _7I4731_$1I4488_$1I4620_DIA;
 reg [1:16] _7I4731_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_159_7 (_7I4731_$1I4488_$1I4620_DIA[7], _7I4731_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_159_6 (_7I4731_$1I4488_$1I4620_DIA[6], _7I4731_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_159_5 (_7I4731_$1I4488_$1I4620_DIA[5], _7I4731_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_159_4 (_7I4731_$1I4488_$1I4620_DIA[4], _7I4731_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_159_3 (_7I4731_$1I4488_$1I4620_DIA[3], _7I4731_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_159_2 (_7I4731_$1I4488_$1I4620_DIA[2], _7I4731_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_159_1 (_7I4731_$1I4488_$1I4620_DIA[1], _7I4731_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_159_0 (_7I4731_$1I4488_$1I4620_DIA[0], _7I4731_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _7I4731_$1I4488_$1I4620_DIB;
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_160_15 (_7I4731_$1I4488_$1I4620_DIB[15], _7I4731_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_160_14 (_7I4731_$1I4488_$1I4620_DIB[14], _7I4731_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_160_13 (_7I4731_$1I4488_$1I4620_DIB[13], _7I4731_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_160_12 (_7I4731_$1I4488_$1I4620_DIB[12], _7I4731_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_160_11 (_7I4731_$1I4488_$1I4620_DIB[11], _7I4731_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_160_10 (_7I4731_$1I4488_$1I4620_DIB[10], _7I4731_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_160_9 (_7I4731_$1I4488_$1I4620_DIB[9], _7I4731_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_160_8 (_7I4731_$1I4488_$1I4620_DIB[8], _7I4731_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_160_7 (_7I4731_$1I4488_$1I4620_DIB[7], _7I4731_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_160_6 (_7I4731_$1I4488_$1I4620_DIB[6], _7I4731_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_160_5 (_7I4731_$1I4488_$1I4620_DIB[5], _7I4731_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_160_4 (_7I4731_$1I4488_$1I4620_DIB[4], _7I4731_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_160_3 (_7I4731_$1I4488_$1I4620_DIB[3], _7I4731_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_160_2 (_7I4731_$1I4488_$1I4620_DIB[2], _7I4731_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_160_1 (_7I4731_$1I4488_$1I4620_DIB[1], _7I4731_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_160_0 (_7I4731_$1I4488_$1I4620_DIB[0], _7I4731_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _7I4731_$1I4488_$1I4620_DIPA;
 reg [1:16] _7I4731_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_161_0 (_7I4731_$1I4488_$1I4620_DIPA[0], _7I4731_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _7I4731_$1I4488_$1I4620_DIPB;
 reg [1:16] _7I4731_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_162_1 (_7I4731_$1I4488_$1I4620_DIPB[1], _7I4731_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _7I4731_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_162_0 (_7I4731_$1I4488_$1I4620_DIPB[0], _7I4731_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _7I4731_$1I4488_$1I4620_ENA;
 reg [1:16] _7I4731_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_163 (_7I4731_$1I4488_$1I4620_ENA, _7I4731_$1I4488_$1I4620_ENA__vlIN);

 wire  _7I4731_$1I4488_$1I4620_ENB;
 reg [1:16] _7I4731_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_164 (_7I4731_$1I4488_$1I4620_ENB, _7I4731_$1I4488_$1I4620_ENB__vlIN);

 wire  _7I4731_$1I4488_$1I4620_SSRA;
 reg [1:16] _7I4731_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_165 (_7I4731_$1I4488_$1I4620_SSRA, _7I4731_$1I4488_$1I4620_SSRA__vlIN);

 wire  _7I4731_$1I4488_$1I4620_SSRB;
 reg [1:16] _7I4731_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_166 (_7I4731_$1I4488_$1I4620_SSRB, _7I4731_$1I4488_$1I4620_SSRB__vlIN);

 wire  _7I4731_$1I4488_$1I4620_WEA;
 reg [1:16] _7I4731_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_167 (_7I4731_$1I4488_$1I4620_WEA, _7I4731_$1I4488_$1I4620_WEA__vlIN);

 wire  _7I4731_$1I4488_$1I4620_WEB;
 reg [1:16] _7I4731_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_168 (_7I4731_$1I4488_$1I4620_WEB, _7I4731_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _7I4731_$1I4488_$1I4620 ( _7I4731_$1I4488_$1I4620_DOA , _7I4731_$1I4488_$1I4620_DOB , _7I4731_$1I4488_$1I4620_DOPA , _7I4731_$1I4488_$1I4620_DOPB , _7I4731_$1I4488_$1I4620_ADDRA , _7I4731_$1I4488_$1I4620_ADDRB , _7I4731_$1I4488_$1I4620_CLKA , _7I4731_$1I4488_$1I4620_CLKB , _7I4731_$1I4488_$1I4620_DIA , _7I4731_$1I4488_$1I4620_DIB , _7I4731_$1I4488_$1I4620_DIPA , _7I4731_$1I4488_$1I4620_DIPB , _7I4731_$1I4488_$1I4620_ENA , _7I4731_$1I4488_$1I4620_ENB , _7I4731_$1I4488_$1I4620_SSRA , _7I4731_$1I4488_$1I4620_SSRB , _7I4731_$1I4488_$1I4620_WEA , _7I4731_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4712_$1I4488_$1I4621_DOA;

 wire [15:0] _7I4712_$1I4488_$1I4621_DOB;

 wire [0:0] _7I4712_$1I4488_$1I4621_DOPA;

 wire [1:0] _7I4712_$1I4488_$1I4621_DOPB;

 wire [10:0] _7I4712_$1I4488_$1I4621_ADDRA;
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_169_10 (_7I4712_$1I4488_$1I4621_ADDRA[10], _7I4712_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_169_9 (_7I4712_$1I4488_$1I4621_ADDRA[9], _7I4712_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_169_8 (_7I4712_$1I4488_$1I4621_ADDRA[8], _7I4712_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_169_7 (_7I4712_$1I4488_$1I4621_ADDRA[7], _7I4712_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_169_6 (_7I4712_$1I4488_$1I4621_ADDRA[6], _7I4712_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_169_5 (_7I4712_$1I4488_$1I4621_ADDRA[5], _7I4712_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_169_4 (_7I4712_$1I4488_$1I4621_ADDRA[4], _7I4712_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_169_3 (_7I4712_$1I4488_$1I4621_ADDRA[3], _7I4712_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_169_2 (_7I4712_$1I4488_$1I4621_ADDRA[2], _7I4712_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_169_1 (_7I4712_$1I4488_$1I4621_ADDRA[1], _7I4712_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_169_0 (_7I4712_$1I4488_$1I4621_ADDRA[0], _7I4712_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _7I4712_$1I4488_$1I4621_ADDRB;
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_170_9 (_7I4712_$1I4488_$1I4621_ADDRB[9], _7I4712_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_170_8 (_7I4712_$1I4488_$1I4621_ADDRB[8], _7I4712_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_170_7 (_7I4712_$1I4488_$1I4621_ADDRB[7], _7I4712_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_170_6 (_7I4712_$1I4488_$1I4621_ADDRB[6], _7I4712_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_170_5 (_7I4712_$1I4488_$1I4621_ADDRB[5], _7I4712_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_170_4 (_7I4712_$1I4488_$1I4621_ADDRB[4], _7I4712_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_170_3 (_7I4712_$1I4488_$1I4621_ADDRB[3], _7I4712_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_170_2 (_7I4712_$1I4488_$1I4621_ADDRB[2], _7I4712_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_170_1 (_7I4712_$1I4488_$1I4621_ADDRB[1], _7I4712_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_170_0 (_7I4712_$1I4488_$1I4621_ADDRB[0], _7I4712_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _7I4712_$1I4488_$1I4621_CLKA;
 reg [1:16] _7I4712_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_171 (_7I4712_$1I4488_$1I4621_CLKA, _7I4712_$1I4488_$1I4621_CLKA__vlIN);

 wire  _7I4712_$1I4488_$1I4621_CLKB;
 reg [1:16] _7I4712_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_172 (_7I4712_$1I4488_$1I4621_CLKB, _7I4712_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _7I4712_$1I4488_$1I4621_DIA;
 reg [1:16] _7I4712_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_173_7 (_7I4712_$1I4488_$1I4621_DIA[7], _7I4712_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_173_6 (_7I4712_$1I4488_$1I4621_DIA[6], _7I4712_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_173_5 (_7I4712_$1I4488_$1I4621_DIA[5], _7I4712_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_173_4 (_7I4712_$1I4488_$1I4621_DIA[4], _7I4712_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_173_3 (_7I4712_$1I4488_$1I4621_DIA[3], _7I4712_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_173_2 (_7I4712_$1I4488_$1I4621_DIA[2], _7I4712_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_173_1 (_7I4712_$1I4488_$1I4621_DIA[1], _7I4712_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_173_0 (_7I4712_$1I4488_$1I4621_DIA[0], _7I4712_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _7I4712_$1I4488_$1I4621_DIB;
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_174_15 (_7I4712_$1I4488_$1I4621_DIB[15], _7I4712_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_174_14 (_7I4712_$1I4488_$1I4621_DIB[14], _7I4712_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_174_13 (_7I4712_$1I4488_$1I4621_DIB[13], _7I4712_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_174_12 (_7I4712_$1I4488_$1I4621_DIB[12], _7I4712_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_174_11 (_7I4712_$1I4488_$1I4621_DIB[11], _7I4712_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_174_10 (_7I4712_$1I4488_$1I4621_DIB[10], _7I4712_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_174_9 (_7I4712_$1I4488_$1I4621_DIB[9], _7I4712_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_174_8 (_7I4712_$1I4488_$1I4621_DIB[8], _7I4712_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_174_7 (_7I4712_$1I4488_$1I4621_DIB[7], _7I4712_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_174_6 (_7I4712_$1I4488_$1I4621_DIB[6], _7I4712_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_174_5 (_7I4712_$1I4488_$1I4621_DIB[5], _7I4712_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_174_4 (_7I4712_$1I4488_$1I4621_DIB[4], _7I4712_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_174_3 (_7I4712_$1I4488_$1I4621_DIB[3], _7I4712_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_174_2 (_7I4712_$1I4488_$1I4621_DIB[2], _7I4712_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_174_1 (_7I4712_$1I4488_$1I4621_DIB[1], _7I4712_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_174_0 (_7I4712_$1I4488_$1I4621_DIB[0], _7I4712_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _7I4712_$1I4488_$1I4621_DIPA;
 reg [1:16] _7I4712_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_175_0 (_7I4712_$1I4488_$1I4621_DIPA[0], _7I4712_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _7I4712_$1I4488_$1I4621_DIPB;
 reg [1:16] _7I4712_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_176_1 (_7I4712_$1I4488_$1I4621_DIPB[1], _7I4712_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_176_0 (_7I4712_$1I4488_$1I4621_DIPB[0], _7I4712_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _7I4712_$1I4488_$1I4621_ENA;
 reg [1:16] _7I4712_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_177 (_7I4712_$1I4488_$1I4621_ENA, _7I4712_$1I4488_$1I4621_ENA__vlIN);

 wire  _7I4712_$1I4488_$1I4621_ENB;
 reg [1:16] _7I4712_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_178 (_7I4712_$1I4488_$1I4621_ENB, _7I4712_$1I4488_$1I4621_ENB__vlIN);

 wire  _7I4712_$1I4488_$1I4621_SSRA;
 reg [1:16] _7I4712_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_179 (_7I4712_$1I4488_$1I4621_SSRA, _7I4712_$1I4488_$1I4621_SSRA__vlIN);

 wire  _7I4712_$1I4488_$1I4621_SSRB;
 reg [1:16] _7I4712_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_180 (_7I4712_$1I4488_$1I4621_SSRB, _7I4712_$1I4488_$1I4621_SSRB__vlIN);

 wire  _7I4712_$1I4488_$1I4621_WEA;
 reg [1:16] _7I4712_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_181 (_7I4712_$1I4488_$1I4621_WEA, _7I4712_$1I4488_$1I4621_WEA__vlIN);

 wire  _7I4712_$1I4488_$1I4621_WEB;
 reg [1:16] _7I4712_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_182 (_7I4712_$1I4488_$1I4621_WEB, _7I4712_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _7I4712_$1I4488_$1I4621 ( _7I4712_$1I4488_$1I4621_DOA , _7I4712_$1I4488_$1I4621_DOB , _7I4712_$1I4488_$1I4621_DOPA , _7I4712_$1I4488_$1I4621_DOPB , _7I4712_$1I4488_$1I4621_ADDRA , _7I4712_$1I4488_$1I4621_ADDRB , _7I4712_$1I4488_$1I4621_CLKA , _7I4712_$1I4488_$1I4621_CLKB , _7I4712_$1I4488_$1I4621_DIA , _7I4712_$1I4488_$1I4621_DIB , _7I4712_$1I4488_$1I4621_DIPA , _7I4712_$1I4488_$1I4621_DIPB , _7I4712_$1I4488_$1I4621_ENA , _7I4712_$1I4488_$1I4621_ENB , _7I4712_$1I4488_$1I4621_SSRA , _7I4712_$1I4488_$1I4621_SSRB , _7I4712_$1I4488_$1I4621_WEA , _7I4712_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4712_$1I4488_$1I4620_DOA;

 wire [15:0] _7I4712_$1I4488_$1I4620_DOB;

 wire [0:0] _7I4712_$1I4488_$1I4620_DOPA;

 wire [1:0] _7I4712_$1I4488_$1I4620_DOPB;

 wire [10:0] _7I4712_$1I4488_$1I4620_ADDRA;
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_183_10 (_7I4712_$1I4488_$1I4620_ADDRA[10], _7I4712_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_183_9 (_7I4712_$1I4488_$1I4620_ADDRA[9], _7I4712_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_183_8 (_7I4712_$1I4488_$1I4620_ADDRA[8], _7I4712_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_183_7 (_7I4712_$1I4488_$1I4620_ADDRA[7], _7I4712_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_183_6 (_7I4712_$1I4488_$1I4620_ADDRA[6], _7I4712_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_183_5 (_7I4712_$1I4488_$1I4620_ADDRA[5], _7I4712_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_183_4 (_7I4712_$1I4488_$1I4620_ADDRA[4], _7I4712_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_183_3 (_7I4712_$1I4488_$1I4620_ADDRA[3], _7I4712_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_183_2 (_7I4712_$1I4488_$1I4620_ADDRA[2], _7I4712_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_183_1 (_7I4712_$1I4488_$1I4620_ADDRA[1], _7I4712_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_183_0 (_7I4712_$1I4488_$1I4620_ADDRA[0], _7I4712_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _7I4712_$1I4488_$1I4620_ADDRB;
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_184_9 (_7I4712_$1I4488_$1I4620_ADDRB[9], _7I4712_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_184_8 (_7I4712_$1I4488_$1I4620_ADDRB[8], _7I4712_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_184_7 (_7I4712_$1I4488_$1I4620_ADDRB[7], _7I4712_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_184_6 (_7I4712_$1I4488_$1I4620_ADDRB[6], _7I4712_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_184_5 (_7I4712_$1I4488_$1I4620_ADDRB[5], _7I4712_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_184_4 (_7I4712_$1I4488_$1I4620_ADDRB[4], _7I4712_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_184_3 (_7I4712_$1I4488_$1I4620_ADDRB[3], _7I4712_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_184_2 (_7I4712_$1I4488_$1I4620_ADDRB[2], _7I4712_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_184_1 (_7I4712_$1I4488_$1I4620_ADDRB[1], _7I4712_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_184_0 (_7I4712_$1I4488_$1I4620_ADDRB[0], _7I4712_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _7I4712_$1I4488_$1I4620_CLKA;
 reg [1:16] _7I4712_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_185 (_7I4712_$1I4488_$1I4620_CLKA, _7I4712_$1I4488_$1I4620_CLKA__vlIN);

 wire  _7I4712_$1I4488_$1I4620_CLKB;
 reg [1:16] _7I4712_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_186 (_7I4712_$1I4488_$1I4620_CLKB, _7I4712_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _7I4712_$1I4488_$1I4620_DIA;
 reg [1:16] _7I4712_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_187_7 (_7I4712_$1I4488_$1I4620_DIA[7], _7I4712_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_187_6 (_7I4712_$1I4488_$1I4620_DIA[6], _7I4712_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_187_5 (_7I4712_$1I4488_$1I4620_DIA[5], _7I4712_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_187_4 (_7I4712_$1I4488_$1I4620_DIA[4], _7I4712_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_187_3 (_7I4712_$1I4488_$1I4620_DIA[3], _7I4712_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_187_2 (_7I4712_$1I4488_$1I4620_DIA[2], _7I4712_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_187_1 (_7I4712_$1I4488_$1I4620_DIA[1], _7I4712_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_187_0 (_7I4712_$1I4488_$1I4620_DIA[0], _7I4712_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _7I4712_$1I4488_$1I4620_DIB;
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_188_15 (_7I4712_$1I4488_$1I4620_DIB[15], _7I4712_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_188_14 (_7I4712_$1I4488_$1I4620_DIB[14], _7I4712_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_188_13 (_7I4712_$1I4488_$1I4620_DIB[13], _7I4712_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_188_12 (_7I4712_$1I4488_$1I4620_DIB[12], _7I4712_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_188_11 (_7I4712_$1I4488_$1I4620_DIB[11], _7I4712_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_188_10 (_7I4712_$1I4488_$1I4620_DIB[10], _7I4712_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_188_9 (_7I4712_$1I4488_$1I4620_DIB[9], _7I4712_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_188_8 (_7I4712_$1I4488_$1I4620_DIB[8], _7I4712_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_188_7 (_7I4712_$1I4488_$1I4620_DIB[7], _7I4712_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_188_6 (_7I4712_$1I4488_$1I4620_DIB[6], _7I4712_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_188_5 (_7I4712_$1I4488_$1I4620_DIB[5], _7I4712_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_188_4 (_7I4712_$1I4488_$1I4620_DIB[4], _7I4712_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_188_3 (_7I4712_$1I4488_$1I4620_DIB[3], _7I4712_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_188_2 (_7I4712_$1I4488_$1I4620_DIB[2], _7I4712_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_188_1 (_7I4712_$1I4488_$1I4620_DIB[1], _7I4712_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_188_0 (_7I4712_$1I4488_$1I4620_DIB[0], _7I4712_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _7I4712_$1I4488_$1I4620_DIPA;
 reg [1:16] _7I4712_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_189_0 (_7I4712_$1I4488_$1I4620_DIPA[0], _7I4712_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _7I4712_$1I4488_$1I4620_DIPB;
 reg [1:16] _7I4712_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_190_1 (_7I4712_$1I4488_$1I4620_DIPB[1], _7I4712_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _7I4712_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_190_0 (_7I4712_$1I4488_$1I4620_DIPB[0], _7I4712_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _7I4712_$1I4488_$1I4620_ENA;
 reg [1:16] _7I4712_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_191 (_7I4712_$1I4488_$1I4620_ENA, _7I4712_$1I4488_$1I4620_ENA__vlIN);

 wire  _7I4712_$1I4488_$1I4620_ENB;
 reg [1:16] _7I4712_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_192 (_7I4712_$1I4488_$1I4620_ENB, _7I4712_$1I4488_$1I4620_ENB__vlIN);

 wire  _7I4712_$1I4488_$1I4620_SSRA;
 reg [1:16] _7I4712_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_193 (_7I4712_$1I4488_$1I4620_SSRA, _7I4712_$1I4488_$1I4620_SSRA__vlIN);

 wire  _7I4712_$1I4488_$1I4620_SSRB;
 reg [1:16] _7I4712_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_194 (_7I4712_$1I4488_$1I4620_SSRB, _7I4712_$1I4488_$1I4620_SSRB__vlIN);

 wire  _7I4712_$1I4488_$1I4620_WEA;
 reg [1:16] _7I4712_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_195 (_7I4712_$1I4488_$1I4620_WEA, _7I4712_$1I4488_$1I4620_WEA__vlIN);

 wire  _7I4712_$1I4488_$1I4620_WEB;
 reg [1:16] _7I4712_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_196 (_7I4712_$1I4488_$1I4620_WEB, _7I4712_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _7I4712_$1I4488_$1I4620 ( _7I4712_$1I4488_$1I4620_DOA , _7I4712_$1I4488_$1I4620_DOB , _7I4712_$1I4488_$1I4620_DOPA , _7I4712_$1I4488_$1I4620_DOPB , _7I4712_$1I4488_$1I4620_ADDRA , _7I4712_$1I4488_$1I4620_ADDRB , _7I4712_$1I4488_$1I4620_CLKA , _7I4712_$1I4488_$1I4620_CLKB , _7I4712_$1I4488_$1I4620_DIA , _7I4712_$1I4488_$1I4620_DIB , _7I4712_$1I4488_$1I4620_DIPA , _7I4712_$1I4488_$1I4620_DIPB , _7I4712_$1I4488_$1I4620_ENA , _7I4712_$1I4488_$1I4620_ENB , _7I4712_$1I4488_$1I4620_SSRA , _7I4712_$1I4488_$1I4620_SSRB , _7I4712_$1I4488_$1I4620_WEA , _7I4712_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4651_$1I4488_$1I4621_DOA;

 wire [15:0] _7I4651_$1I4488_$1I4621_DOB;

 wire [0:0] _7I4651_$1I4488_$1I4621_DOPA;

 wire [1:0] _7I4651_$1I4488_$1I4621_DOPB;

 wire [10:0] _7I4651_$1I4488_$1I4621_ADDRA;
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_197_10 (_7I4651_$1I4488_$1I4621_ADDRA[10], _7I4651_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_197_9 (_7I4651_$1I4488_$1I4621_ADDRA[9], _7I4651_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_197_8 (_7I4651_$1I4488_$1I4621_ADDRA[8], _7I4651_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_197_7 (_7I4651_$1I4488_$1I4621_ADDRA[7], _7I4651_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_197_6 (_7I4651_$1I4488_$1I4621_ADDRA[6], _7I4651_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_197_5 (_7I4651_$1I4488_$1I4621_ADDRA[5], _7I4651_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_197_4 (_7I4651_$1I4488_$1I4621_ADDRA[4], _7I4651_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_197_3 (_7I4651_$1I4488_$1I4621_ADDRA[3], _7I4651_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_197_2 (_7I4651_$1I4488_$1I4621_ADDRA[2], _7I4651_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_197_1 (_7I4651_$1I4488_$1I4621_ADDRA[1], _7I4651_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_197_0 (_7I4651_$1I4488_$1I4621_ADDRA[0], _7I4651_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _7I4651_$1I4488_$1I4621_ADDRB;
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_198_9 (_7I4651_$1I4488_$1I4621_ADDRB[9], _7I4651_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_198_8 (_7I4651_$1I4488_$1I4621_ADDRB[8], _7I4651_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_198_7 (_7I4651_$1I4488_$1I4621_ADDRB[7], _7I4651_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_198_6 (_7I4651_$1I4488_$1I4621_ADDRB[6], _7I4651_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_198_5 (_7I4651_$1I4488_$1I4621_ADDRB[5], _7I4651_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_198_4 (_7I4651_$1I4488_$1I4621_ADDRB[4], _7I4651_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_198_3 (_7I4651_$1I4488_$1I4621_ADDRB[3], _7I4651_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_198_2 (_7I4651_$1I4488_$1I4621_ADDRB[2], _7I4651_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_198_1 (_7I4651_$1I4488_$1I4621_ADDRB[1], _7I4651_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_198_0 (_7I4651_$1I4488_$1I4621_ADDRB[0], _7I4651_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _7I4651_$1I4488_$1I4621_CLKA;
 reg [1:16] _7I4651_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_199 (_7I4651_$1I4488_$1I4621_CLKA, _7I4651_$1I4488_$1I4621_CLKA__vlIN);

 wire  _7I4651_$1I4488_$1I4621_CLKB;
 reg [1:16] _7I4651_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_200 (_7I4651_$1I4488_$1I4621_CLKB, _7I4651_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _7I4651_$1I4488_$1I4621_DIA;
 reg [1:16] _7I4651_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_201_7 (_7I4651_$1I4488_$1I4621_DIA[7], _7I4651_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_201_6 (_7I4651_$1I4488_$1I4621_DIA[6], _7I4651_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_201_5 (_7I4651_$1I4488_$1I4621_DIA[5], _7I4651_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_201_4 (_7I4651_$1I4488_$1I4621_DIA[4], _7I4651_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_201_3 (_7I4651_$1I4488_$1I4621_DIA[3], _7I4651_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_201_2 (_7I4651_$1I4488_$1I4621_DIA[2], _7I4651_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_201_1 (_7I4651_$1I4488_$1I4621_DIA[1], _7I4651_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_201_0 (_7I4651_$1I4488_$1I4621_DIA[0], _7I4651_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _7I4651_$1I4488_$1I4621_DIB;
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_202_15 (_7I4651_$1I4488_$1I4621_DIB[15], _7I4651_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_202_14 (_7I4651_$1I4488_$1I4621_DIB[14], _7I4651_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_202_13 (_7I4651_$1I4488_$1I4621_DIB[13], _7I4651_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_202_12 (_7I4651_$1I4488_$1I4621_DIB[12], _7I4651_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_202_11 (_7I4651_$1I4488_$1I4621_DIB[11], _7I4651_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_202_10 (_7I4651_$1I4488_$1I4621_DIB[10], _7I4651_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_202_9 (_7I4651_$1I4488_$1I4621_DIB[9], _7I4651_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_202_8 (_7I4651_$1I4488_$1I4621_DIB[8], _7I4651_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_202_7 (_7I4651_$1I4488_$1I4621_DIB[7], _7I4651_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_202_6 (_7I4651_$1I4488_$1I4621_DIB[6], _7I4651_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_202_5 (_7I4651_$1I4488_$1I4621_DIB[5], _7I4651_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_202_4 (_7I4651_$1I4488_$1I4621_DIB[4], _7I4651_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_202_3 (_7I4651_$1I4488_$1I4621_DIB[3], _7I4651_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_202_2 (_7I4651_$1I4488_$1I4621_DIB[2], _7I4651_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_202_1 (_7I4651_$1I4488_$1I4621_DIB[1], _7I4651_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_202_0 (_7I4651_$1I4488_$1I4621_DIB[0], _7I4651_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _7I4651_$1I4488_$1I4621_DIPA;
 reg [1:16] _7I4651_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_203_0 (_7I4651_$1I4488_$1I4621_DIPA[0], _7I4651_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _7I4651_$1I4488_$1I4621_DIPB;
 reg [1:16] _7I4651_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_204_1 (_7I4651_$1I4488_$1I4621_DIPB[1], _7I4651_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_204_0 (_7I4651_$1I4488_$1I4621_DIPB[0], _7I4651_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _7I4651_$1I4488_$1I4621_ENA;
 reg [1:16] _7I4651_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_205 (_7I4651_$1I4488_$1I4621_ENA, _7I4651_$1I4488_$1I4621_ENA__vlIN);

 wire  _7I4651_$1I4488_$1I4621_ENB;
 reg [1:16] _7I4651_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_206 (_7I4651_$1I4488_$1I4621_ENB, _7I4651_$1I4488_$1I4621_ENB__vlIN);

 wire  _7I4651_$1I4488_$1I4621_SSRA;
 reg [1:16] _7I4651_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_207 (_7I4651_$1I4488_$1I4621_SSRA, _7I4651_$1I4488_$1I4621_SSRA__vlIN);

 wire  _7I4651_$1I4488_$1I4621_SSRB;
 reg [1:16] _7I4651_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_208 (_7I4651_$1I4488_$1I4621_SSRB, _7I4651_$1I4488_$1I4621_SSRB__vlIN);

 wire  _7I4651_$1I4488_$1I4621_WEA;
 reg [1:16] _7I4651_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_209 (_7I4651_$1I4488_$1I4621_WEA, _7I4651_$1I4488_$1I4621_WEA__vlIN);

 wire  _7I4651_$1I4488_$1I4621_WEB;
 reg [1:16] _7I4651_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_210 (_7I4651_$1I4488_$1I4621_WEB, _7I4651_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _7I4651_$1I4488_$1I4621 ( _7I4651_$1I4488_$1I4621_DOA , _7I4651_$1I4488_$1I4621_DOB , _7I4651_$1I4488_$1I4621_DOPA , _7I4651_$1I4488_$1I4621_DOPB , _7I4651_$1I4488_$1I4621_ADDRA , _7I4651_$1I4488_$1I4621_ADDRB , _7I4651_$1I4488_$1I4621_CLKA , _7I4651_$1I4488_$1I4621_CLKB , _7I4651_$1I4488_$1I4621_DIA , _7I4651_$1I4488_$1I4621_DIB , _7I4651_$1I4488_$1I4621_DIPA , _7I4651_$1I4488_$1I4621_DIPB , _7I4651_$1I4488_$1I4621_ENA , _7I4651_$1I4488_$1I4621_ENB , _7I4651_$1I4488_$1I4621_SSRA , _7I4651_$1I4488_$1I4621_SSRB , _7I4651_$1I4488_$1I4621_WEA , _7I4651_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4651_$1I4488_$1I4620_DOA;

 wire [15:0] _7I4651_$1I4488_$1I4620_DOB;

 wire [0:0] _7I4651_$1I4488_$1I4620_DOPA;

 wire [1:0] _7I4651_$1I4488_$1I4620_DOPB;

 wire [10:0] _7I4651_$1I4488_$1I4620_ADDRA;
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_211_10 (_7I4651_$1I4488_$1I4620_ADDRA[10], _7I4651_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_211_9 (_7I4651_$1I4488_$1I4620_ADDRA[9], _7I4651_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_211_8 (_7I4651_$1I4488_$1I4620_ADDRA[8], _7I4651_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_211_7 (_7I4651_$1I4488_$1I4620_ADDRA[7], _7I4651_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_211_6 (_7I4651_$1I4488_$1I4620_ADDRA[6], _7I4651_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_211_5 (_7I4651_$1I4488_$1I4620_ADDRA[5], _7I4651_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_211_4 (_7I4651_$1I4488_$1I4620_ADDRA[4], _7I4651_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_211_3 (_7I4651_$1I4488_$1I4620_ADDRA[3], _7I4651_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_211_2 (_7I4651_$1I4488_$1I4620_ADDRA[2], _7I4651_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_211_1 (_7I4651_$1I4488_$1I4620_ADDRA[1], _7I4651_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_211_0 (_7I4651_$1I4488_$1I4620_ADDRA[0], _7I4651_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _7I4651_$1I4488_$1I4620_ADDRB;
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_212_9 (_7I4651_$1I4488_$1I4620_ADDRB[9], _7I4651_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_212_8 (_7I4651_$1I4488_$1I4620_ADDRB[8], _7I4651_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_212_7 (_7I4651_$1I4488_$1I4620_ADDRB[7], _7I4651_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_212_6 (_7I4651_$1I4488_$1I4620_ADDRB[6], _7I4651_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_212_5 (_7I4651_$1I4488_$1I4620_ADDRB[5], _7I4651_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_212_4 (_7I4651_$1I4488_$1I4620_ADDRB[4], _7I4651_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_212_3 (_7I4651_$1I4488_$1I4620_ADDRB[3], _7I4651_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_212_2 (_7I4651_$1I4488_$1I4620_ADDRB[2], _7I4651_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_212_1 (_7I4651_$1I4488_$1I4620_ADDRB[1], _7I4651_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_212_0 (_7I4651_$1I4488_$1I4620_ADDRB[0], _7I4651_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _7I4651_$1I4488_$1I4620_CLKA;
 reg [1:16] _7I4651_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_213 (_7I4651_$1I4488_$1I4620_CLKA, _7I4651_$1I4488_$1I4620_CLKA__vlIN);

 wire  _7I4651_$1I4488_$1I4620_CLKB;
 reg [1:16] _7I4651_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_214 (_7I4651_$1I4488_$1I4620_CLKB, _7I4651_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _7I4651_$1I4488_$1I4620_DIA;
 reg [1:16] _7I4651_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_215_7 (_7I4651_$1I4488_$1I4620_DIA[7], _7I4651_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_215_6 (_7I4651_$1I4488_$1I4620_DIA[6], _7I4651_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_215_5 (_7I4651_$1I4488_$1I4620_DIA[5], _7I4651_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_215_4 (_7I4651_$1I4488_$1I4620_DIA[4], _7I4651_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_215_3 (_7I4651_$1I4488_$1I4620_DIA[3], _7I4651_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_215_2 (_7I4651_$1I4488_$1I4620_DIA[2], _7I4651_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_215_1 (_7I4651_$1I4488_$1I4620_DIA[1], _7I4651_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_215_0 (_7I4651_$1I4488_$1I4620_DIA[0], _7I4651_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _7I4651_$1I4488_$1I4620_DIB;
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_216_15 (_7I4651_$1I4488_$1I4620_DIB[15], _7I4651_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_216_14 (_7I4651_$1I4488_$1I4620_DIB[14], _7I4651_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_216_13 (_7I4651_$1I4488_$1I4620_DIB[13], _7I4651_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_216_12 (_7I4651_$1I4488_$1I4620_DIB[12], _7I4651_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_216_11 (_7I4651_$1I4488_$1I4620_DIB[11], _7I4651_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_216_10 (_7I4651_$1I4488_$1I4620_DIB[10], _7I4651_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_216_9 (_7I4651_$1I4488_$1I4620_DIB[9], _7I4651_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_216_8 (_7I4651_$1I4488_$1I4620_DIB[8], _7I4651_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_216_7 (_7I4651_$1I4488_$1I4620_DIB[7], _7I4651_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_216_6 (_7I4651_$1I4488_$1I4620_DIB[6], _7I4651_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_216_5 (_7I4651_$1I4488_$1I4620_DIB[5], _7I4651_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_216_4 (_7I4651_$1I4488_$1I4620_DIB[4], _7I4651_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_216_3 (_7I4651_$1I4488_$1I4620_DIB[3], _7I4651_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_216_2 (_7I4651_$1I4488_$1I4620_DIB[2], _7I4651_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_216_1 (_7I4651_$1I4488_$1I4620_DIB[1], _7I4651_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_216_0 (_7I4651_$1I4488_$1I4620_DIB[0], _7I4651_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _7I4651_$1I4488_$1I4620_DIPA;
 reg [1:16] _7I4651_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_217_0 (_7I4651_$1I4488_$1I4620_DIPA[0], _7I4651_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _7I4651_$1I4488_$1I4620_DIPB;
 reg [1:16] _7I4651_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_218_1 (_7I4651_$1I4488_$1I4620_DIPB[1], _7I4651_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _7I4651_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_218_0 (_7I4651_$1I4488_$1I4620_DIPB[0], _7I4651_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _7I4651_$1I4488_$1I4620_ENA;
 reg [1:16] _7I4651_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_219 (_7I4651_$1I4488_$1I4620_ENA, _7I4651_$1I4488_$1I4620_ENA__vlIN);

 wire  _7I4651_$1I4488_$1I4620_ENB;
 reg [1:16] _7I4651_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_220 (_7I4651_$1I4488_$1I4620_ENB, _7I4651_$1I4488_$1I4620_ENB__vlIN);

 wire  _7I4651_$1I4488_$1I4620_SSRA;
 reg [1:16] _7I4651_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_221 (_7I4651_$1I4488_$1I4620_SSRA, _7I4651_$1I4488_$1I4620_SSRA__vlIN);

 wire  _7I4651_$1I4488_$1I4620_SSRB;
 reg [1:16] _7I4651_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_222 (_7I4651_$1I4488_$1I4620_SSRB, _7I4651_$1I4488_$1I4620_SSRB__vlIN);

 wire  _7I4651_$1I4488_$1I4620_WEA;
 reg [1:16] _7I4651_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_223 (_7I4651_$1I4488_$1I4620_WEA, _7I4651_$1I4488_$1I4620_WEA__vlIN);

 wire  _7I4651_$1I4488_$1I4620_WEB;
 reg [1:16] _7I4651_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_224 (_7I4651_$1I4488_$1I4620_WEB, _7I4651_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _7I4651_$1I4488_$1I4620 ( _7I4651_$1I4488_$1I4620_DOA , _7I4651_$1I4488_$1I4620_DOB , _7I4651_$1I4488_$1I4620_DOPA , _7I4651_$1I4488_$1I4620_DOPB , _7I4651_$1I4488_$1I4620_ADDRA , _7I4651_$1I4488_$1I4620_ADDRB , _7I4651_$1I4488_$1I4620_CLKA , _7I4651_$1I4488_$1I4620_CLKB , _7I4651_$1I4488_$1I4620_DIA , _7I4651_$1I4488_$1I4620_DIB , _7I4651_$1I4488_$1I4620_DIPA , _7I4651_$1I4488_$1I4620_DIPB , _7I4651_$1I4488_$1I4620_ENA , _7I4651_$1I4488_$1I4620_ENB , _7I4651_$1I4488_$1I4620_SSRA , _7I4651_$1I4488_$1I4620_SSRB , _7I4651_$1I4488_$1I4620_WEA , _7I4651_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4632_$1I4488_$1I4621_DOA;

 wire [15:0] _7I4632_$1I4488_$1I4621_DOB;

 wire [0:0] _7I4632_$1I4488_$1I4621_DOPA;

 wire [1:0] _7I4632_$1I4488_$1I4621_DOPB;

 wire [10:0] _7I4632_$1I4488_$1I4621_ADDRA;
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_225_10 (_7I4632_$1I4488_$1I4621_ADDRA[10], _7I4632_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_225_9 (_7I4632_$1I4488_$1I4621_ADDRA[9], _7I4632_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_225_8 (_7I4632_$1I4488_$1I4621_ADDRA[8], _7I4632_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_225_7 (_7I4632_$1I4488_$1I4621_ADDRA[7], _7I4632_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_225_6 (_7I4632_$1I4488_$1I4621_ADDRA[6], _7I4632_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_225_5 (_7I4632_$1I4488_$1I4621_ADDRA[5], _7I4632_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_225_4 (_7I4632_$1I4488_$1I4621_ADDRA[4], _7I4632_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_225_3 (_7I4632_$1I4488_$1I4621_ADDRA[3], _7I4632_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_225_2 (_7I4632_$1I4488_$1I4621_ADDRA[2], _7I4632_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_225_1 (_7I4632_$1I4488_$1I4621_ADDRA[1], _7I4632_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_225_0 (_7I4632_$1I4488_$1I4621_ADDRA[0], _7I4632_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _7I4632_$1I4488_$1I4621_ADDRB;
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_226_9 (_7I4632_$1I4488_$1I4621_ADDRB[9], _7I4632_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_226_8 (_7I4632_$1I4488_$1I4621_ADDRB[8], _7I4632_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_226_7 (_7I4632_$1I4488_$1I4621_ADDRB[7], _7I4632_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_226_6 (_7I4632_$1I4488_$1I4621_ADDRB[6], _7I4632_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_226_5 (_7I4632_$1I4488_$1I4621_ADDRB[5], _7I4632_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_226_4 (_7I4632_$1I4488_$1I4621_ADDRB[4], _7I4632_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_226_3 (_7I4632_$1I4488_$1I4621_ADDRB[3], _7I4632_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_226_2 (_7I4632_$1I4488_$1I4621_ADDRB[2], _7I4632_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_226_1 (_7I4632_$1I4488_$1I4621_ADDRB[1], _7I4632_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_226_0 (_7I4632_$1I4488_$1I4621_ADDRB[0], _7I4632_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _7I4632_$1I4488_$1I4621_CLKA;
 reg [1:16] _7I4632_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_227 (_7I4632_$1I4488_$1I4621_CLKA, _7I4632_$1I4488_$1I4621_CLKA__vlIN);

 wire  _7I4632_$1I4488_$1I4621_CLKB;
 reg [1:16] _7I4632_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_228 (_7I4632_$1I4488_$1I4621_CLKB, _7I4632_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _7I4632_$1I4488_$1I4621_DIA;
 reg [1:16] _7I4632_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_229_7 (_7I4632_$1I4488_$1I4621_DIA[7], _7I4632_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_229_6 (_7I4632_$1I4488_$1I4621_DIA[6], _7I4632_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_229_5 (_7I4632_$1I4488_$1I4621_DIA[5], _7I4632_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_229_4 (_7I4632_$1I4488_$1I4621_DIA[4], _7I4632_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_229_3 (_7I4632_$1I4488_$1I4621_DIA[3], _7I4632_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_229_2 (_7I4632_$1I4488_$1I4621_DIA[2], _7I4632_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_229_1 (_7I4632_$1I4488_$1I4621_DIA[1], _7I4632_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_229_0 (_7I4632_$1I4488_$1I4621_DIA[0], _7I4632_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _7I4632_$1I4488_$1I4621_DIB;
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_230_15 (_7I4632_$1I4488_$1I4621_DIB[15], _7I4632_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_230_14 (_7I4632_$1I4488_$1I4621_DIB[14], _7I4632_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_230_13 (_7I4632_$1I4488_$1I4621_DIB[13], _7I4632_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_230_12 (_7I4632_$1I4488_$1I4621_DIB[12], _7I4632_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_230_11 (_7I4632_$1I4488_$1I4621_DIB[11], _7I4632_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_230_10 (_7I4632_$1I4488_$1I4621_DIB[10], _7I4632_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_230_9 (_7I4632_$1I4488_$1I4621_DIB[9], _7I4632_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_230_8 (_7I4632_$1I4488_$1I4621_DIB[8], _7I4632_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_230_7 (_7I4632_$1I4488_$1I4621_DIB[7], _7I4632_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_230_6 (_7I4632_$1I4488_$1I4621_DIB[6], _7I4632_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_230_5 (_7I4632_$1I4488_$1I4621_DIB[5], _7I4632_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_230_4 (_7I4632_$1I4488_$1I4621_DIB[4], _7I4632_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_230_3 (_7I4632_$1I4488_$1I4621_DIB[3], _7I4632_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_230_2 (_7I4632_$1I4488_$1I4621_DIB[2], _7I4632_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_230_1 (_7I4632_$1I4488_$1I4621_DIB[1], _7I4632_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_230_0 (_7I4632_$1I4488_$1I4621_DIB[0], _7I4632_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _7I4632_$1I4488_$1I4621_DIPA;
 reg [1:16] _7I4632_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_231_0 (_7I4632_$1I4488_$1I4621_DIPA[0], _7I4632_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _7I4632_$1I4488_$1I4621_DIPB;
 reg [1:16] _7I4632_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_232_1 (_7I4632_$1I4488_$1I4621_DIPB[1], _7I4632_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_232_0 (_7I4632_$1I4488_$1I4621_DIPB[0], _7I4632_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _7I4632_$1I4488_$1I4621_ENA;
 reg [1:16] _7I4632_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_233 (_7I4632_$1I4488_$1I4621_ENA, _7I4632_$1I4488_$1I4621_ENA__vlIN);

 wire  _7I4632_$1I4488_$1I4621_ENB;
 reg [1:16] _7I4632_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_234 (_7I4632_$1I4488_$1I4621_ENB, _7I4632_$1I4488_$1I4621_ENB__vlIN);

 wire  _7I4632_$1I4488_$1I4621_SSRA;
 reg [1:16] _7I4632_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_235 (_7I4632_$1I4488_$1I4621_SSRA, _7I4632_$1I4488_$1I4621_SSRA__vlIN);

 wire  _7I4632_$1I4488_$1I4621_SSRB;
 reg [1:16] _7I4632_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_236 (_7I4632_$1I4488_$1I4621_SSRB, _7I4632_$1I4488_$1I4621_SSRB__vlIN);

 wire  _7I4632_$1I4488_$1I4621_WEA;
 reg [1:16] _7I4632_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_237 (_7I4632_$1I4488_$1I4621_WEA, _7I4632_$1I4488_$1I4621_WEA__vlIN);

 wire  _7I4632_$1I4488_$1I4621_WEB;
 reg [1:16] _7I4632_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_238 (_7I4632_$1I4488_$1I4621_WEB, _7I4632_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _7I4632_$1I4488_$1I4621 ( _7I4632_$1I4488_$1I4621_DOA , _7I4632_$1I4488_$1I4621_DOB , _7I4632_$1I4488_$1I4621_DOPA , _7I4632_$1I4488_$1I4621_DOPB , _7I4632_$1I4488_$1I4621_ADDRA , _7I4632_$1I4488_$1I4621_ADDRB , _7I4632_$1I4488_$1I4621_CLKA , _7I4632_$1I4488_$1I4621_CLKB , _7I4632_$1I4488_$1I4621_DIA , _7I4632_$1I4488_$1I4621_DIB , _7I4632_$1I4488_$1I4621_DIPA , _7I4632_$1I4488_$1I4621_DIPB , _7I4632_$1I4488_$1I4621_ENA , _7I4632_$1I4488_$1I4621_ENB , _7I4632_$1I4488_$1I4621_SSRA , _7I4632_$1I4488_$1I4621_SSRB , _7I4632_$1I4488_$1I4621_WEA , _7I4632_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4632_$1I4488_$1I4620_DOA;

 wire [15:0] _7I4632_$1I4488_$1I4620_DOB;

 wire [0:0] _7I4632_$1I4488_$1I4620_DOPA;

 wire [1:0] _7I4632_$1I4488_$1I4620_DOPB;

 wire [10:0] _7I4632_$1I4488_$1I4620_ADDRA;
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_239_10 (_7I4632_$1I4488_$1I4620_ADDRA[10], _7I4632_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_239_9 (_7I4632_$1I4488_$1I4620_ADDRA[9], _7I4632_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_239_8 (_7I4632_$1I4488_$1I4620_ADDRA[8], _7I4632_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_239_7 (_7I4632_$1I4488_$1I4620_ADDRA[7], _7I4632_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_239_6 (_7I4632_$1I4488_$1I4620_ADDRA[6], _7I4632_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_239_5 (_7I4632_$1I4488_$1I4620_ADDRA[5], _7I4632_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_239_4 (_7I4632_$1I4488_$1I4620_ADDRA[4], _7I4632_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_239_3 (_7I4632_$1I4488_$1I4620_ADDRA[3], _7I4632_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_239_2 (_7I4632_$1I4488_$1I4620_ADDRA[2], _7I4632_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_239_1 (_7I4632_$1I4488_$1I4620_ADDRA[1], _7I4632_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_239_0 (_7I4632_$1I4488_$1I4620_ADDRA[0], _7I4632_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _7I4632_$1I4488_$1I4620_ADDRB;
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_240_9 (_7I4632_$1I4488_$1I4620_ADDRB[9], _7I4632_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_240_8 (_7I4632_$1I4488_$1I4620_ADDRB[8], _7I4632_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_240_7 (_7I4632_$1I4488_$1I4620_ADDRB[7], _7I4632_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_240_6 (_7I4632_$1I4488_$1I4620_ADDRB[6], _7I4632_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_240_5 (_7I4632_$1I4488_$1I4620_ADDRB[5], _7I4632_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_240_4 (_7I4632_$1I4488_$1I4620_ADDRB[4], _7I4632_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_240_3 (_7I4632_$1I4488_$1I4620_ADDRB[3], _7I4632_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_240_2 (_7I4632_$1I4488_$1I4620_ADDRB[2], _7I4632_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_240_1 (_7I4632_$1I4488_$1I4620_ADDRB[1], _7I4632_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_240_0 (_7I4632_$1I4488_$1I4620_ADDRB[0], _7I4632_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _7I4632_$1I4488_$1I4620_CLKA;
 reg [1:16] _7I4632_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_241 (_7I4632_$1I4488_$1I4620_CLKA, _7I4632_$1I4488_$1I4620_CLKA__vlIN);

 wire  _7I4632_$1I4488_$1I4620_CLKB;
 reg [1:16] _7I4632_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_242 (_7I4632_$1I4488_$1I4620_CLKB, _7I4632_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _7I4632_$1I4488_$1I4620_DIA;
 reg [1:16] _7I4632_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_243_7 (_7I4632_$1I4488_$1I4620_DIA[7], _7I4632_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_243_6 (_7I4632_$1I4488_$1I4620_DIA[6], _7I4632_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_243_5 (_7I4632_$1I4488_$1I4620_DIA[5], _7I4632_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_243_4 (_7I4632_$1I4488_$1I4620_DIA[4], _7I4632_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_243_3 (_7I4632_$1I4488_$1I4620_DIA[3], _7I4632_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_243_2 (_7I4632_$1I4488_$1I4620_DIA[2], _7I4632_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_243_1 (_7I4632_$1I4488_$1I4620_DIA[1], _7I4632_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_243_0 (_7I4632_$1I4488_$1I4620_DIA[0], _7I4632_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _7I4632_$1I4488_$1I4620_DIB;
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_244_15 (_7I4632_$1I4488_$1I4620_DIB[15], _7I4632_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_244_14 (_7I4632_$1I4488_$1I4620_DIB[14], _7I4632_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_244_13 (_7I4632_$1I4488_$1I4620_DIB[13], _7I4632_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_244_12 (_7I4632_$1I4488_$1I4620_DIB[12], _7I4632_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_244_11 (_7I4632_$1I4488_$1I4620_DIB[11], _7I4632_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_244_10 (_7I4632_$1I4488_$1I4620_DIB[10], _7I4632_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_244_9 (_7I4632_$1I4488_$1I4620_DIB[9], _7I4632_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_244_8 (_7I4632_$1I4488_$1I4620_DIB[8], _7I4632_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_244_7 (_7I4632_$1I4488_$1I4620_DIB[7], _7I4632_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_244_6 (_7I4632_$1I4488_$1I4620_DIB[6], _7I4632_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_244_5 (_7I4632_$1I4488_$1I4620_DIB[5], _7I4632_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_244_4 (_7I4632_$1I4488_$1I4620_DIB[4], _7I4632_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_244_3 (_7I4632_$1I4488_$1I4620_DIB[3], _7I4632_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_244_2 (_7I4632_$1I4488_$1I4620_DIB[2], _7I4632_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_244_1 (_7I4632_$1I4488_$1I4620_DIB[1], _7I4632_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_244_0 (_7I4632_$1I4488_$1I4620_DIB[0], _7I4632_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _7I4632_$1I4488_$1I4620_DIPA;
 reg [1:16] _7I4632_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_245_0 (_7I4632_$1I4488_$1I4620_DIPA[0], _7I4632_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _7I4632_$1I4488_$1I4620_DIPB;
 reg [1:16] _7I4632_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_246_1 (_7I4632_$1I4488_$1I4620_DIPB[1], _7I4632_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _7I4632_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_246_0 (_7I4632_$1I4488_$1I4620_DIPB[0], _7I4632_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _7I4632_$1I4488_$1I4620_ENA;
 reg [1:16] _7I4632_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_247 (_7I4632_$1I4488_$1I4620_ENA, _7I4632_$1I4488_$1I4620_ENA__vlIN);

 wire  _7I4632_$1I4488_$1I4620_ENB;
 reg [1:16] _7I4632_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_248 (_7I4632_$1I4488_$1I4620_ENB, _7I4632_$1I4488_$1I4620_ENB__vlIN);

 wire  _7I4632_$1I4488_$1I4620_SSRA;
 reg [1:16] _7I4632_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_249 (_7I4632_$1I4488_$1I4620_SSRA, _7I4632_$1I4488_$1I4620_SSRA__vlIN);

 wire  _7I4632_$1I4488_$1I4620_SSRB;
 reg [1:16] _7I4632_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_250 (_7I4632_$1I4488_$1I4620_SSRB, _7I4632_$1I4488_$1I4620_SSRB__vlIN);

 wire  _7I4632_$1I4488_$1I4620_WEA;
 reg [1:16] _7I4632_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_251 (_7I4632_$1I4488_$1I4620_WEA, _7I4632_$1I4488_$1I4620_WEA__vlIN);

 wire  _7I4632_$1I4488_$1I4620_WEB;
 reg [1:16] _7I4632_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_252 (_7I4632_$1I4488_$1I4620_WEB, _7I4632_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _7I4632_$1I4488_$1I4620 ( _7I4632_$1I4488_$1I4620_DOA , _7I4632_$1I4488_$1I4620_DOB , _7I4632_$1I4488_$1I4620_DOPA , _7I4632_$1I4488_$1I4620_DOPB , _7I4632_$1I4488_$1I4620_ADDRA , _7I4632_$1I4488_$1I4620_ADDRB , _7I4632_$1I4488_$1I4620_CLKA , _7I4632_$1I4488_$1I4620_CLKB , _7I4632_$1I4488_$1I4620_DIA , _7I4632_$1I4488_$1I4620_DIB , _7I4632_$1I4488_$1I4620_DIPA , _7I4632_$1I4488_$1I4620_DIPB , _7I4632_$1I4488_$1I4620_ENA , _7I4632_$1I4488_$1I4620_ENB , _7I4632_$1I4488_$1I4620_SSRA , _7I4632_$1I4488_$1I4620_SSRB , _7I4632_$1I4488_$1I4620_WEA , _7I4632_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4616_$1I4488_$1I4621_DOA;

 wire [15:0] _7I4616_$1I4488_$1I4621_DOB;

 wire [0:0] _7I4616_$1I4488_$1I4621_DOPA;

 wire [1:0] _7I4616_$1I4488_$1I4621_DOPB;

 wire [10:0] _7I4616_$1I4488_$1I4621_ADDRA;
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_253_10 (_7I4616_$1I4488_$1I4621_ADDRA[10], _7I4616_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_253_9 (_7I4616_$1I4488_$1I4621_ADDRA[9], _7I4616_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_253_8 (_7I4616_$1I4488_$1I4621_ADDRA[8], _7I4616_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_253_7 (_7I4616_$1I4488_$1I4621_ADDRA[7], _7I4616_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_253_6 (_7I4616_$1I4488_$1I4621_ADDRA[6], _7I4616_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_253_5 (_7I4616_$1I4488_$1I4621_ADDRA[5], _7I4616_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_253_4 (_7I4616_$1I4488_$1I4621_ADDRA[4], _7I4616_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_253_3 (_7I4616_$1I4488_$1I4621_ADDRA[3], _7I4616_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_253_2 (_7I4616_$1I4488_$1I4621_ADDRA[2], _7I4616_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_253_1 (_7I4616_$1I4488_$1I4621_ADDRA[1], _7I4616_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_253_0 (_7I4616_$1I4488_$1I4621_ADDRA[0], _7I4616_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _7I4616_$1I4488_$1I4621_ADDRB;
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_254_9 (_7I4616_$1I4488_$1I4621_ADDRB[9], _7I4616_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_254_8 (_7I4616_$1I4488_$1I4621_ADDRB[8], _7I4616_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_254_7 (_7I4616_$1I4488_$1I4621_ADDRB[7], _7I4616_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_254_6 (_7I4616_$1I4488_$1I4621_ADDRB[6], _7I4616_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_254_5 (_7I4616_$1I4488_$1I4621_ADDRB[5], _7I4616_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_254_4 (_7I4616_$1I4488_$1I4621_ADDRB[4], _7I4616_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_254_3 (_7I4616_$1I4488_$1I4621_ADDRB[3], _7I4616_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_254_2 (_7I4616_$1I4488_$1I4621_ADDRB[2], _7I4616_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_254_1 (_7I4616_$1I4488_$1I4621_ADDRB[1], _7I4616_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_254_0 (_7I4616_$1I4488_$1I4621_ADDRB[0], _7I4616_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _7I4616_$1I4488_$1I4621_CLKA;
 reg [1:16] _7I4616_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_255 (_7I4616_$1I4488_$1I4621_CLKA, _7I4616_$1I4488_$1I4621_CLKA__vlIN);

 wire  _7I4616_$1I4488_$1I4621_CLKB;
 reg [1:16] _7I4616_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_256 (_7I4616_$1I4488_$1I4621_CLKB, _7I4616_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _7I4616_$1I4488_$1I4621_DIA;
 reg [1:16] _7I4616_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_257_7 (_7I4616_$1I4488_$1I4621_DIA[7], _7I4616_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_257_6 (_7I4616_$1I4488_$1I4621_DIA[6], _7I4616_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_257_5 (_7I4616_$1I4488_$1I4621_DIA[5], _7I4616_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_257_4 (_7I4616_$1I4488_$1I4621_DIA[4], _7I4616_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_257_3 (_7I4616_$1I4488_$1I4621_DIA[3], _7I4616_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_257_2 (_7I4616_$1I4488_$1I4621_DIA[2], _7I4616_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_257_1 (_7I4616_$1I4488_$1I4621_DIA[1], _7I4616_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_257_0 (_7I4616_$1I4488_$1I4621_DIA[0], _7I4616_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _7I4616_$1I4488_$1I4621_DIB;
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_258_15 (_7I4616_$1I4488_$1I4621_DIB[15], _7I4616_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_258_14 (_7I4616_$1I4488_$1I4621_DIB[14], _7I4616_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_258_13 (_7I4616_$1I4488_$1I4621_DIB[13], _7I4616_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_258_12 (_7I4616_$1I4488_$1I4621_DIB[12], _7I4616_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_258_11 (_7I4616_$1I4488_$1I4621_DIB[11], _7I4616_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_258_10 (_7I4616_$1I4488_$1I4621_DIB[10], _7I4616_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_258_9 (_7I4616_$1I4488_$1I4621_DIB[9], _7I4616_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_258_8 (_7I4616_$1I4488_$1I4621_DIB[8], _7I4616_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_258_7 (_7I4616_$1I4488_$1I4621_DIB[7], _7I4616_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_258_6 (_7I4616_$1I4488_$1I4621_DIB[6], _7I4616_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_258_5 (_7I4616_$1I4488_$1I4621_DIB[5], _7I4616_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_258_4 (_7I4616_$1I4488_$1I4621_DIB[4], _7I4616_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_258_3 (_7I4616_$1I4488_$1I4621_DIB[3], _7I4616_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_258_2 (_7I4616_$1I4488_$1I4621_DIB[2], _7I4616_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_258_1 (_7I4616_$1I4488_$1I4621_DIB[1], _7I4616_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_258_0 (_7I4616_$1I4488_$1I4621_DIB[0], _7I4616_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _7I4616_$1I4488_$1I4621_DIPA;
 reg [1:16] _7I4616_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_259_0 (_7I4616_$1I4488_$1I4621_DIPA[0], _7I4616_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _7I4616_$1I4488_$1I4621_DIPB;
 reg [1:16] _7I4616_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_260_1 (_7I4616_$1I4488_$1I4621_DIPB[1], _7I4616_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_260_0 (_7I4616_$1I4488_$1I4621_DIPB[0], _7I4616_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _7I4616_$1I4488_$1I4621_ENA;
 reg [1:16] _7I4616_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_261 (_7I4616_$1I4488_$1I4621_ENA, _7I4616_$1I4488_$1I4621_ENA__vlIN);

 wire  _7I4616_$1I4488_$1I4621_ENB;
 reg [1:16] _7I4616_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_262 (_7I4616_$1I4488_$1I4621_ENB, _7I4616_$1I4488_$1I4621_ENB__vlIN);

 wire  _7I4616_$1I4488_$1I4621_SSRA;
 reg [1:16] _7I4616_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_263 (_7I4616_$1I4488_$1I4621_SSRA, _7I4616_$1I4488_$1I4621_SSRA__vlIN);

 wire  _7I4616_$1I4488_$1I4621_SSRB;
 reg [1:16] _7I4616_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_264 (_7I4616_$1I4488_$1I4621_SSRB, _7I4616_$1I4488_$1I4621_SSRB__vlIN);

 wire  _7I4616_$1I4488_$1I4621_WEA;
 reg [1:16] _7I4616_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_265 (_7I4616_$1I4488_$1I4621_WEA, _7I4616_$1I4488_$1I4621_WEA__vlIN);

 wire  _7I4616_$1I4488_$1I4621_WEB;
 reg [1:16] _7I4616_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_266 (_7I4616_$1I4488_$1I4621_WEB, _7I4616_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _7I4616_$1I4488_$1I4621 ( _7I4616_$1I4488_$1I4621_DOA , _7I4616_$1I4488_$1I4621_DOB , _7I4616_$1I4488_$1I4621_DOPA , _7I4616_$1I4488_$1I4621_DOPB , _7I4616_$1I4488_$1I4621_ADDRA , _7I4616_$1I4488_$1I4621_ADDRB , _7I4616_$1I4488_$1I4621_CLKA , _7I4616_$1I4488_$1I4621_CLKB , _7I4616_$1I4488_$1I4621_DIA , _7I4616_$1I4488_$1I4621_DIB , _7I4616_$1I4488_$1I4621_DIPA , _7I4616_$1I4488_$1I4621_DIPB , _7I4616_$1I4488_$1I4621_ENA , _7I4616_$1I4488_$1I4621_ENB , _7I4616_$1I4488_$1I4621_SSRA , _7I4616_$1I4488_$1I4621_SSRB , _7I4616_$1I4488_$1I4621_WEA , _7I4616_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4616_$1I4488_$1I4620_DOA;

 wire [15:0] _7I4616_$1I4488_$1I4620_DOB;

 wire [0:0] _7I4616_$1I4488_$1I4620_DOPA;

 wire [1:0] _7I4616_$1I4488_$1I4620_DOPB;

 wire [10:0] _7I4616_$1I4488_$1I4620_ADDRA;
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_267_10 (_7I4616_$1I4488_$1I4620_ADDRA[10], _7I4616_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_267_9 (_7I4616_$1I4488_$1I4620_ADDRA[9], _7I4616_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_267_8 (_7I4616_$1I4488_$1I4620_ADDRA[8], _7I4616_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_267_7 (_7I4616_$1I4488_$1I4620_ADDRA[7], _7I4616_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_267_6 (_7I4616_$1I4488_$1I4620_ADDRA[6], _7I4616_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_267_5 (_7I4616_$1I4488_$1I4620_ADDRA[5], _7I4616_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_267_4 (_7I4616_$1I4488_$1I4620_ADDRA[4], _7I4616_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_267_3 (_7I4616_$1I4488_$1I4620_ADDRA[3], _7I4616_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_267_2 (_7I4616_$1I4488_$1I4620_ADDRA[2], _7I4616_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_267_1 (_7I4616_$1I4488_$1I4620_ADDRA[1], _7I4616_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_267_0 (_7I4616_$1I4488_$1I4620_ADDRA[0], _7I4616_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _7I4616_$1I4488_$1I4620_ADDRB;
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_268_9 (_7I4616_$1I4488_$1I4620_ADDRB[9], _7I4616_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_268_8 (_7I4616_$1I4488_$1I4620_ADDRB[8], _7I4616_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_268_7 (_7I4616_$1I4488_$1I4620_ADDRB[7], _7I4616_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_268_6 (_7I4616_$1I4488_$1I4620_ADDRB[6], _7I4616_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_268_5 (_7I4616_$1I4488_$1I4620_ADDRB[5], _7I4616_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_268_4 (_7I4616_$1I4488_$1I4620_ADDRB[4], _7I4616_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_268_3 (_7I4616_$1I4488_$1I4620_ADDRB[3], _7I4616_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_268_2 (_7I4616_$1I4488_$1I4620_ADDRB[2], _7I4616_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_268_1 (_7I4616_$1I4488_$1I4620_ADDRB[1], _7I4616_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_268_0 (_7I4616_$1I4488_$1I4620_ADDRB[0], _7I4616_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _7I4616_$1I4488_$1I4620_CLKA;
 reg [1:16] _7I4616_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_269 (_7I4616_$1I4488_$1I4620_CLKA, _7I4616_$1I4488_$1I4620_CLKA__vlIN);

 wire  _7I4616_$1I4488_$1I4620_CLKB;
 reg [1:16] _7I4616_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_270 (_7I4616_$1I4488_$1I4620_CLKB, _7I4616_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _7I4616_$1I4488_$1I4620_DIA;
 reg [1:16] _7I4616_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_271_7 (_7I4616_$1I4488_$1I4620_DIA[7], _7I4616_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_271_6 (_7I4616_$1I4488_$1I4620_DIA[6], _7I4616_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_271_5 (_7I4616_$1I4488_$1I4620_DIA[5], _7I4616_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_271_4 (_7I4616_$1I4488_$1I4620_DIA[4], _7I4616_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_271_3 (_7I4616_$1I4488_$1I4620_DIA[3], _7I4616_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_271_2 (_7I4616_$1I4488_$1I4620_DIA[2], _7I4616_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_271_1 (_7I4616_$1I4488_$1I4620_DIA[1], _7I4616_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_271_0 (_7I4616_$1I4488_$1I4620_DIA[0], _7I4616_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _7I4616_$1I4488_$1I4620_DIB;
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_272_15 (_7I4616_$1I4488_$1I4620_DIB[15], _7I4616_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_272_14 (_7I4616_$1I4488_$1I4620_DIB[14], _7I4616_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_272_13 (_7I4616_$1I4488_$1I4620_DIB[13], _7I4616_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_272_12 (_7I4616_$1I4488_$1I4620_DIB[12], _7I4616_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_272_11 (_7I4616_$1I4488_$1I4620_DIB[11], _7I4616_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_272_10 (_7I4616_$1I4488_$1I4620_DIB[10], _7I4616_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_272_9 (_7I4616_$1I4488_$1I4620_DIB[9], _7I4616_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_272_8 (_7I4616_$1I4488_$1I4620_DIB[8], _7I4616_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_272_7 (_7I4616_$1I4488_$1I4620_DIB[7], _7I4616_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_272_6 (_7I4616_$1I4488_$1I4620_DIB[6], _7I4616_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_272_5 (_7I4616_$1I4488_$1I4620_DIB[5], _7I4616_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_272_4 (_7I4616_$1I4488_$1I4620_DIB[4], _7I4616_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_272_3 (_7I4616_$1I4488_$1I4620_DIB[3], _7I4616_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_272_2 (_7I4616_$1I4488_$1I4620_DIB[2], _7I4616_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_272_1 (_7I4616_$1I4488_$1I4620_DIB[1], _7I4616_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_272_0 (_7I4616_$1I4488_$1I4620_DIB[0], _7I4616_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _7I4616_$1I4488_$1I4620_DIPA;
 reg [1:16] _7I4616_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_273_0 (_7I4616_$1I4488_$1I4620_DIPA[0], _7I4616_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _7I4616_$1I4488_$1I4620_DIPB;
 reg [1:16] _7I4616_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_274_1 (_7I4616_$1I4488_$1I4620_DIPB[1], _7I4616_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _7I4616_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_274_0 (_7I4616_$1I4488_$1I4620_DIPB[0], _7I4616_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _7I4616_$1I4488_$1I4620_ENA;
 reg [1:16] _7I4616_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_275 (_7I4616_$1I4488_$1I4620_ENA, _7I4616_$1I4488_$1I4620_ENA__vlIN);

 wire  _7I4616_$1I4488_$1I4620_ENB;
 reg [1:16] _7I4616_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_276 (_7I4616_$1I4488_$1I4620_ENB, _7I4616_$1I4488_$1I4620_ENB__vlIN);

 wire  _7I4616_$1I4488_$1I4620_SSRA;
 reg [1:16] _7I4616_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_277 (_7I4616_$1I4488_$1I4620_SSRA, _7I4616_$1I4488_$1I4620_SSRA__vlIN);

 wire  _7I4616_$1I4488_$1I4620_SSRB;
 reg [1:16] _7I4616_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_278 (_7I4616_$1I4488_$1I4620_SSRB, _7I4616_$1I4488_$1I4620_SSRB__vlIN);

 wire  _7I4616_$1I4488_$1I4620_WEA;
 reg [1:16] _7I4616_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_279 (_7I4616_$1I4488_$1I4620_WEA, _7I4616_$1I4488_$1I4620_WEA__vlIN);

 wire  _7I4616_$1I4488_$1I4620_WEB;
 reg [1:16] _7I4616_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_280 (_7I4616_$1I4488_$1I4620_WEB, _7I4616_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _7I4616_$1I4488_$1I4620 ( _7I4616_$1I4488_$1I4620_DOA , _7I4616_$1I4488_$1I4620_DOB , _7I4616_$1I4488_$1I4620_DOPA , _7I4616_$1I4488_$1I4620_DOPB , _7I4616_$1I4488_$1I4620_ADDRA , _7I4616_$1I4488_$1I4620_ADDRB , _7I4616_$1I4488_$1I4620_CLKA , _7I4616_$1I4488_$1I4620_CLKB , _7I4616_$1I4488_$1I4620_DIA , _7I4616_$1I4488_$1I4620_DIB , _7I4616_$1I4488_$1I4620_DIPA , _7I4616_$1I4488_$1I4620_DIPB , _7I4616_$1I4488_$1I4620_ENA , _7I4616_$1I4488_$1I4620_ENB , _7I4616_$1I4488_$1I4620_SSRA , _7I4616_$1I4488_$1I4620_SSRB , _7I4616_$1I4488_$1I4620_WEA , _7I4616_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4615_$1I4488_$1I4621_DOA;

 wire [15:0] _7I4615_$1I4488_$1I4621_DOB;

 wire [0:0] _7I4615_$1I4488_$1I4621_DOPA;

 wire [1:0] _7I4615_$1I4488_$1I4621_DOPB;

 wire [10:0] _7I4615_$1I4488_$1I4621_ADDRA;
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_281_10 (_7I4615_$1I4488_$1I4621_ADDRA[10], _7I4615_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_281_9 (_7I4615_$1I4488_$1I4621_ADDRA[9], _7I4615_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_281_8 (_7I4615_$1I4488_$1I4621_ADDRA[8], _7I4615_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_281_7 (_7I4615_$1I4488_$1I4621_ADDRA[7], _7I4615_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_281_6 (_7I4615_$1I4488_$1I4621_ADDRA[6], _7I4615_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_281_5 (_7I4615_$1I4488_$1I4621_ADDRA[5], _7I4615_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_281_4 (_7I4615_$1I4488_$1I4621_ADDRA[4], _7I4615_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_281_3 (_7I4615_$1I4488_$1I4621_ADDRA[3], _7I4615_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_281_2 (_7I4615_$1I4488_$1I4621_ADDRA[2], _7I4615_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_281_1 (_7I4615_$1I4488_$1I4621_ADDRA[1], _7I4615_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_281_0 (_7I4615_$1I4488_$1I4621_ADDRA[0], _7I4615_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _7I4615_$1I4488_$1I4621_ADDRB;
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_282_9 (_7I4615_$1I4488_$1I4621_ADDRB[9], _7I4615_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_282_8 (_7I4615_$1I4488_$1I4621_ADDRB[8], _7I4615_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_282_7 (_7I4615_$1I4488_$1I4621_ADDRB[7], _7I4615_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_282_6 (_7I4615_$1I4488_$1I4621_ADDRB[6], _7I4615_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_282_5 (_7I4615_$1I4488_$1I4621_ADDRB[5], _7I4615_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_282_4 (_7I4615_$1I4488_$1I4621_ADDRB[4], _7I4615_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_282_3 (_7I4615_$1I4488_$1I4621_ADDRB[3], _7I4615_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_282_2 (_7I4615_$1I4488_$1I4621_ADDRB[2], _7I4615_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_282_1 (_7I4615_$1I4488_$1I4621_ADDRB[1], _7I4615_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_282_0 (_7I4615_$1I4488_$1I4621_ADDRB[0], _7I4615_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _7I4615_$1I4488_$1I4621_CLKA;
 reg [1:16] _7I4615_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_283 (_7I4615_$1I4488_$1I4621_CLKA, _7I4615_$1I4488_$1I4621_CLKA__vlIN);

 wire  _7I4615_$1I4488_$1I4621_CLKB;
 reg [1:16] _7I4615_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_284 (_7I4615_$1I4488_$1I4621_CLKB, _7I4615_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _7I4615_$1I4488_$1I4621_DIA;
 reg [1:16] _7I4615_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_285_7 (_7I4615_$1I4488_$1I4621_DIA[7], _7I4615_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_285_6 (_7I4615_$1I4488_$1I4621_DIA[6], _7I4615_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_285_5 (_7I4615_$1I4488_$1I4621_DIA[5], _7I4615_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_285_4 (_7I4615_$1I4488_$1I4621_DIA[4], _7I4615_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_285_3 (_7I4615_$1I4488_$1I4621_DIA[3], _7I4615_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_285_2 (_7I4615_$1I4488_$1I4621_DIA[2], _7I4615_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_285_1 (_7I4615_$1I4488_$1I4621_DIA[1], _7I4615_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_285_0 (_7I4615_$1I4488_$1I4621_DIA[0], _7I4615_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _7I4615_$1I4488_$1I4621_DIB;
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_286_15 (_7I4615_$1I4488_$1I4621_DIB[15], _7I4615_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_286_14 (_7I4615_$1I4488_$1I4621_DIB[14], _7I4615_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_286_13 (_7I4615_$1I4488_$1I4621_DIB[13], _7I4615_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_286_12 (_7I4615_$1I4488_$1I4621_DIB[12], _7I4615_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_286_11 (_7I4615_$1I4488_$1I4621_DIB[11], _7I4615_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_286_10 (_7I4615_$1I4488_$1I4621_DIB[10], _7I4615_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_286_9 (_7I4615_$1I4488_$1I4621_DIB[9], _7I4615_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_286_8 (_7I4615_$1I4488_$1I4621_DIB[8], _7I4615_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_286_7 (_7I4615_$1I4488_$1I4621_DIB[7], _7I4615_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_286_6 (_7I4615_$1I4488_$1I4621_DIB[6], _7I4615_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_286_5 (_7I4615_$1I4488_$1I4621_DIB[5], _7I4615_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_286_4 (_7I4615_$1I4488_$1I4621_DIB[4], _7I4615_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_286_3 (_7I4615_$1I4488_$1I4621_DIB[3], _7I4615_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_286_2 (_7I4615_$1I4488_$1I4621_DIB[2], _7I4615_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_286_1 (_7I4615_$1I4488_$1I4621_DIB[1], _7I4615_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_286_0 (_7I4615_$1I4488_$1I4621_DIB[0], _7I4615_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _7I4615_$1I4488_$1I4621_DIPA;
 reg [1:16] _7I4615_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_287_0 (_7I4615_$1I4488_$1I4621_DIPA[0], _7I4615_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _7I4615_$1I4488_$1I4621_DIPB;
 reg [1:16] _7I4615_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_288_1 (_7I4615_$1I4488_$1I4621_DIPB[1], _7I4615_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_288_0 (_7I4615_$1I4488_$1I4621_DIPB[0], _7I4615_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _7I4615_$1I4488_$1I4621_ENA;
 reg [1:16] _7I4615_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_289 (_7I4615_$1I4488_$1I4621_ENA, _7I4615_$1I4488_$1I4621_ENA__vlIN);

 wire  _7I4615_$1I4488_$1I4621_ENB;
 reg [1:16] _7I4615_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_290 (_7I4615_$1I4488_$1I4621_ENB, _7I4615_$1I4488_$1I4621_ENB__vlIN);

 wire  _7I4615_$1I4488_$1I4621_SSRA;
 reg [1:16] _7I4615_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_291 (_7I4615_$1I4488_$1I4621_SSRA, _7I4615_$1I4488_$1I4621_SSRA__vlIN);

 wire  _7I4615_$1I4488_$1I4621_SSRB;
 reg [1:16] _7I4615_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_292 (_7I4615_$1I4488_$1I4621_SSRB, _7I4615_$1I4488_$1I4621_SSRB__vlIN);

 wire  _7I4615_$1I4488_$1I4621_WEA;
 reg [1:16] _7I4615_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_293 (_7I4615_$1I4488_$1I4621_WEA, _7I4615_$1I4488_$1I4621_WEA__vlIN);

 wire  _7I4615_$1I4488_$1I4621_WEB;
 reg [1:16] _7I4615_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_294 (_7I4615_$1I4488_$1I4621_WEB, _7I4615_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _7I4615_$1I4488_$1I4621 ( _7I4615_$1I4488_$1I4621_DOA , _7I4615_$1I4488_$1I4621_DOB , _7I4615_$1I4488_$1I4621_DOPA , _7I4615_$1I4488_$1I4621_DOPB , _7I4615_$1I4488_$1I4621_ADDRA , _7I4615_$1I4488_$1I4621_ADDRB , _7I4615_$1I4488_$1I4621_CLKA , _7I4615_$1I4488_$1I4621_CLKB , _7I4615_$1I4488_$1I4621_DIA , _7I4615_$1I4488_$1I4621_DIB , _7I4615_$1I4488_$1I4621_DIPA , _7I4615_$1I4488_$1I4621_DIPB , _7I4615_$1I4488_$1I4621_ENA , _7I4615_$1I4488_$1I4621_ENB , _7I4615_$1I4488_$1I4621_SSRA , _7I4615_$1I4488_$1I4621_SSRB , _7I4615_$1I4488_$1I4621_WEA , _7I4615_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4615_$1I4488_$1I4620_DOA;

 wire [15:0] _7I4615_$1I4488_$1I4620_DOB;

 wire [0:0] _7I4615_$1I4488_$1I4620_DOPA;

 wire [1:0] _7I4615_$1I4488_$1I4620_DOPB;

 wire [10:0] _7I4615_$1I4488_$1I4620_ADDRA;
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_295_10 (_7I4615_$1I4488_$1I4620_ADDRA[10], _7I4615_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_295_9 (_7I4615_$1I4488_$1I4620_ADDRA[9], _7I4615_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_295_8 (_7I4615_$1I4488_$1I4620_ADDRA[8], _7I4615_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_295_7 (_7I4615_$1I4488_$1I4620_ADDRA[7], _7I4615_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_295_6 (_7I4615_$1I4488_$1I4620_ADDRA[6], _7I4615_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_295_5 (_7I4615_$1I4488_$1I4620_ADDRA[5], _7I4615_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_295_4 (_7I4615_$1I4488_$1I4620_ADDRA[4], _7I4615_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_295_3 (_7I4615_$1I4488_$1I4620_ADDRA[3], _7I4615_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_295_2 (_7I4615_$1I4488_$1I4620_ADDRA[2], _7I4615_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_295_1 (_7I4615_$1I4488_$1I4620_ADDRA[1], _7I4615_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_295_0 (_7I4615_$1I4488_$1I4620_ADDRA[0], _7I4615_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _7I4615_$1I4488_$1I4620_ADDRB;
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_296_9 (_7I4615_$1I4488_$1I4620_ADDRB[9], _7I4615_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_296_8 (_7I4615_$1I4488_$1I4620_ADDRB[8], _7I4615_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_296_7 (_7I4615_$1I4488_$1I4620_ADDRB[7], _7I4615_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_296_6 (_7I4615_$1I4488_$1I4620_ADDRB[6], _7I4615_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_296_5 (_7I4615_$1I4488_$1I4620_ADDRB[5], _7I4615_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_296_4 (_7I4615_$1I4488_$1I4620_ADDRB[4], _7I4615_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_296_3 (_7I4615_$1I4488_$1I4620_ADDRB[3], _7I4615_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_296_2 (_7I4615_$1I4488_$1I4620_ADDRB[2], _7I4615_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_296_1 (_7I4615_$1I4488_$1I4620_ADDRB[1], _7I4615_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_296_0 (_7I4615_$1I4488_$1I4620_ADDRB[0], _7I4615_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _7I4615_$1I4488_$1I4620_CLKA;
 reg [1:16] _7I4615_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_297 (_7I4615_$1I4488_$1I4620_CLKA, _7I4615_$1I4488_$1I4620_CLKA__vlIN);

 wire  _7I4615_$1I4488_$1I4620_CLKB;
 reg [1:16] _7I4615_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_298 (_7I4615_$1I4488_$1I4620_CLKB, _7I4615_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _7I4615_$1I4488_$1I4620_DIA;
 reg [1:16] _7I4615_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_299_7 (_7I4615_$1I4488_$1I4620_DIA[7], _7I4615_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_299_6 (_7I4615_$1I4488_$1I4620_DIA[6], _7I4615_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_299_5 (_7I4615_$1I4488_$1I4620_DIA[5], _7I4615_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_299_4 (_7I4615_$1I4488_$1I4620_DIA[4], _7I4615_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_299_3 (_7I4615_$1I4488_$1I4620_DIA[3], _7I4615_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_299_2 (_7I4615_$1I4488_$1I4620_DIA[2], _7I4615_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_299_1 (_7I4615_$1I4488_$1I4620_DIA[1], _7I4615_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_299_0 (_7I4615_$1I4488_$1I4620_DIA[0], _7I4615_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _7I4615_$1I4488_$1I4620_DIB;
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_300_15 (_7I4615_$1I4488_$1I4620_DIB[15], _7I4615_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_300_14 (_7I4615_$1I4488_$1I4620_DIB[14], _7I4615_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_300_13 (_7I4615_$1I4488_$1I4620_DIB[13], _7I4615_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_300_12 (_7I4615_$1I4488_$1I4620_DIB[12], _7I4615_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_300_11 (_7I4615_$1I4488_$1I4620_DIB[11], _7I4615_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_300_10 (_7I4615_$1I4488_$1I4620_DIB[10], _7I4615_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_300_9 (_7I4615_$1I4488_$1I4620_DIB[9], _7I4615_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_300_8 (_7I4615_$1I4488_$1I4620_DIB[8], _7I4615_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_300_7 (_7I4615_$1I4488_$1I4620_DIB[7], _7I4615_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_300_6 (_7I4615_$1I4488_$1I4620_DIB[6], _7I4615_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_300_5 (_7I4615_$1I4488_$1I4620_DIB[5], _7I4615_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_300_4 (_7I4615_$1I4488_$1I4620_DIB[4], _7I4615_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_300_3 (_7I4615_$1I4488_$1I4620_DIB[3], _7I4615_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_300_2 (_7I4615_$1I4488_$1I4620_DIB[2], _7I4615_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_300_1 (_7I4615_$1I4488_$1I4620_DIB[1], _7I4615_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_300_0 (_7I4615_$1I4488_$1I4620_DIB[0], _7I4615_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _7I4615_$1I4488_$1I4620_DIPA;
 reg [1:16] _7I4615_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_301_0 (_7I4615_$1I4488_$1I4620_DIPA[0], _7I4615_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _7I4615_$1I4488_$1I4620_DIPB;
 reg [1:16] _7I4615_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_302_1 (_7I4615_$1I4488_$1I4620_DIPB[1], _7I4615_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _7I4615_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_302_0 (_7I4615_$1I4488_$1I4620_DIPB[0], _7I4615_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _7I4615_$1I4488_$1I4620_ENA;
 reg [1:16] _7I4615_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_303 (_7I4615_$1I4488_$1I4620_ENA, _7I4615_$1I4488_$1I4620_ENA__vlIN);

 wire  _7I4615_$1I4488_$1I4620_ENB;
 reg [1:16] _7I4615_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_304 (_7I4615_$1I4488_$1I4620_ENB, _7I4615_$1I4488_$1I4620_ENB__vlIN);

 wire  _7I4615_$1I4488_$1I4620_SSRA;
 reg [1:16] _7I4615_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_305 (_7I4615_$1I4488_$1I4620_SSRA, _7I4615_$1I4488_$1I4620_SSRA__vlIN);

 wire  _7I4615_$1I4488_$1I4620_SSRB;
 reg [1:16] _7I4615_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_306 (_7I4615_$1I4488_$1I4620_SSRB, _7I4615_$1I4488_$1I4620_SSRB__vlIN);

 wire  _7I4615_$1I4488_$1I4620_WEA;
 reg [1:16] _7I4615_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_307 (_7I4615_$1I4488_$1I4620_WEA, _7I4615_$1I4488_$1I4620_WEA__vlIN);

 wire  _7I4615_$1I4488_$1I4620_WEB;
 reg [1:16] _7I4615_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_308 (_7I4615_$1I4488_$1I4620_WEB, _7I4615_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _7I4615_$1I4488_$1I4620 ( _7I4615_$1I4488_$1I4620_DOA , _7I4615_$1I4488_$1I4620_DOB , _7I4615_$1I4488_$1I4620_DOPA , _7I4615_$1I4488_$1I4620_DOPB , _7I4615_$1I4488_$1I4620_ADDRA , _7I4615_$1I4488_$1I4620_ADDRB , _7I4615_$1I4488_$1I4620_CLKA , _7I4615_$1I4488_$1I4620_CLKB , _7I4615_$1I4488_$1I4620_DIA , _7I4615_$1I4488_$1I4620_DIB , _7I4615_$1I4488_$1I4620_DIPA , _7I4615_$1I4488_$1I4620_DIPB , _7I4615_$1I4488_$1I4620_ENA , _7I4615_$1I4488_$1I4620_ENB , _7I4615_$1I4488_$1I4620_SSRA , _7I4615_$1I4488_$1I4620_SSRB , _7I4615_$1I4488_$1I4620_WEA , _7I4615_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4614_$1I4488_$1I4621_DOA;

 wire [15:0] _7I4614_$1I4488_$1I4621_DOB;

 wire [0:0] _7I4614_$1I4488_$1I4621_DOPA;

 wire [1:0] _7I4614_$1I4488_$1I4621_DOPB;

 wire [10:0] _7I4614_$1I4488_$1I4621_ADDRA;
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_309_10 (_7I4614_$1I4488_$1I4621_ADDRA[10], _7I4614_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_309_9 (_7I4614_$1I4488_$1I4621_ADDRA[9], _7I4614_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_309_8 (_7I4614_$1I4488_$1I4621_ADDRA[8], _7I4614_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_309_7 (_7I4614_$1I4488_$1I4621_ADDRA[7], _7I4614_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_309_6 (_7I4614_$1I4488_$1I4621_ADDRA[6], _7I4614_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_309_5 (_7I4614_$1I4488_$1I4621_ADDRA[5], _7I4614_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_309_4 (_7I4614_$1I4488_$1I4621_ADDRA[4], _7I4614_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_309_3 (_7I4614_$1I4488_$1I4621_ADDRA[3], _7I4614_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_309_2 (_7I4614_$1I4488_$1I4621_ADDRA[2], _7I4614_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_309_1 (_7I4614_$1I4488_$1I4621_ADDRA[1], _7I4614_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_309_0 (_7I4614_$1I4488_$1I4621_ADDRA[0], _7I4614_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _7I4614_$1I4488_$1I4621_ADDRB;
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_310_9 (_7I4614_$1I4488_$1I4621_ADDRB[9], _7I4614_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_310_8 (_7I4614_$1I4488_$1I4621_ADDRB[8], _7I4614_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_310_7 (_7I4614_$1I4488_$1I4621_ADDRB[7], _7I4614_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_310_6 (_7I4614_$1I4488_$1I4621_ADDRB[6], _7I4614_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_310_5 (_7I4614_$1I4488_$1I4621_ADDRB[5], _7I4614_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_310_4 (_7I4614_$1I4488_$1I4621_ADDRB[4], _7I4614_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_310_3 (_7I4614_$1I4488_$1I4621_ADDRB[3], _7I4614_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_310_2 (_7I4614_$1I4488_$1I4621_ADDRB[2], _7I4614_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_310_1 (_7I4614_$1I4488_$1I4621_ADDRB[1], _7I4614_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_310_0 (_7I4614_$1I4488_$1I4621_ADDRB[0], _7I4614_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _7I4614_$1I4488_$1I4621_CLKA;
 reg [1:16] _7I4614_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_311 (_7I4614_$1I4488_$1I4621_CLKA, _7I4614_$1I4488_$1I4621_CLKA__vlIN);

 wire  _7I4614_$1I4488_$1I4621_CLKB;
 reg [1:16] _7I4614_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_312 (_7I4614_$1I4488_$1I4621_CLKB, _7I4614_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _7I4614_$1I4488_$1I4621_DIA;
 reg [1:16] _7I4614_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_313_7 (_7I4614_$1I4488_$1I4621_DIA[7], _7I4614_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_313_6 (_7I4614_$1I4488_$1I4621_DIA[6], _7I4614_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_313_5 (_7I4614_$1I4488_$1I4621_DIA[5], _7I4614_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_313_4 (_7I4614_$1I4488_$1I4621_DIA[4], _7I4614_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_313_3 (_7I4614_$1I4488_$1I4621_DIA[3], _7I4614_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_313_2 (_7I4614_$1I4488_$1I4621_DIA[2], _7I4614_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_313_1 (_7I4614_$1I4488_$1I4621_DIA[1], _7I4614_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_313_0 (_7I4614_$1I4488_$1I4621_DIA[0], _7I4614_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _7I4614_$1I4488_$1I4621_DIB;
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_314_15 (_7I4614_$1I4488_$1I4621_DIB[15], _7I4614_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_314_14 (_7I4614_$1I4488_$1I4621_DIB[14], _7I4614_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_314_13 (_7I4614_$1I4488_$1I4621_DIB[13], _7I4614_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_314_12 (_7I4614_$1I4488_$1I4621_DIB[12], _7I4614_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_314_11 (_7I4614_$1I4488_$1I4621_DIB[11], _7I4614_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_314_10 (_7I4614_$1I4488_$1I4621_DIB[10], _7I4614_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_314_9 (_7I4614_$1I4488_$1I4621_DIB[9], _7I4614_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_314_8 (_7I4614_$1I4488_$1I4621_DIB[8], _7I4614_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_314_7 (_7I4614_$1I4488_$1I4621_DIB[7], _7I4614_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_314_6 (_7I4614_$1I4488_$1I4621_DIB[6], _7I4614_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_314_5 (_7I4614_$1I4488_$1I4621_DIB[5], _7I4614_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_314_4 (_7I4614_$1I4488_$1I4621_DIB[4], _7I4614_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_314_3 (_7I4614_$1I4488_$1I4621_DIB[3], _7I4614_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_314_2 (_7I4614_$1I4488_$1I4621_DIB[2], _7I4614_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_314_1 (_7I4614_$1I4488_$1I4621_DIB[1], _7I4614_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_314_0 (_7I4614_$1I4488_$1I4621_DIB[0], _7I4614_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _7I4614_$1I4488_$1I4621_DIPA;
 reg [1:16] _7I4614_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_315_0 (_7I4614_$1I4488_$1I4621_DIPA[0], _7I4614_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _7I4614_$1I4488_$1I4621_DIPB;
 reg [1:16] _7I4614_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_316_1 (_7I4614_$1I4488_$1I4621_DIPB[1], _7I4614_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_316_0 (_7I4614_$1I4488_$1I4621_DIPB[0], _7I4614_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _7I4614_$1I4488_$1I4621_ENA;
 reg [1:16] _7I4614_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_317 (_7I4614_$1I4488_$1I4621_ENA, _7I4614_$1I4488_$1I4621_ENA__vlIN);

 wire  _7I4614_$1I4488_$1I4621_ENB;
 reg [1:16] _7I4614_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_318 (_7I4614_$1I4488_$1I4621_ENB, _7I4614_$1I4488_$1I4621_ENB__vlIN);

 wire  _7I4614_$1I4488_$1I4621_SSRA;
 reg [1:16] _7I4614_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_319 (_7I4614_$1I4488_$1I4621_SSRA, _7I4614_$1I4488_$1I4621_SSRA__vlIN);

 wire  _7I4614_$1I4488_$1I4621_SSRB;
 reg [1:16] _7I4614_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_320 (_7I4614_$1I4488_$1I4621_SSRB, _7I4614_$1I4488_$1I4621_SSRB__vlIN);

 wire  _7I4614_$1I4488_$1I4621_WEA;
 reg [1:16] _7I4614_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_321 (_7I4614_$1I4488_$1I4621_WEA, _7I4614_$1I4488_$1I4621_WEA__vlIN);

 wire  _7I4614_$1I4488_$1I4621_WEB;
 reg [1:16] _7I4614_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_322 (_7I4614_$1I4488_$1I4621_WEB, _7I4614_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _7I4614_$1I4488_$1I4621 ( _7I4614_$1I4488_$1I4621_DOA , _7I4614_$1I4488_$1I4621_DOB , _7I4614_$1I4488_$1I4621_DOPA , _7I4614_$1I4488_$1I4621_DOPB , _7I4614_$1I4488_$1I4621_ADDRA , _7I4614_$1I4488_$1I4621_ADDRB , _7I4614_$1I4488_$1I4621_CLKA , _7I4614_$1I4488_$1I4621_CLKB , _7I4614_$1I4488_$1I4621_DIA , _7I4614_$1I4488_$1I4621_DIB , _7I4614_$1I4488_$1I4621_DIPA , _7I4614_$1I4488_$1I4621_DIPB , _7I4614_$1I4488_$1I4621_ENA , _7I4614_$1I4488_$1I4621_ENB , _7I4614_$1I4488_$1I4621_SSRA , _7I4614_$1I4488_$1I4621_SSRB , _7I4614_$1I4488_$1I4621_WEA , _7I4614_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _7I4614_$1I4488_$1I4620_DOA;

 wire [15:0] _7I4614_$1I4488_$1I4620_DOB;

 wire [0:0] _7I4614_$1I4488_$1I4620_DOPA;

 wire [1:0] _7I4614_$1I4488_$1I4620_DOPB;

 wire [10:0] _7I4614_$1I4488_$1I4620_ADDRA;
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_323_10 (_7I4614_$1I4488_$1I4620_ADDRA[10], _7I4614_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_323_9 (_7I4614_$1I4488_$1I4620_ADDRA[9], _7I4614_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_323_8 (_7I4614_$1I4488_$1I4620_ADDRA[8], _7I4614_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_323_7 (_7I4614_$1I4488_$1I4620_ADDRA[7], _7I4614_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_323_6 (_7I4614_$1I4488_$1I4620_ADDRA[6], _7I4614_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_323_5 (_7I4614_$1I4488_$1I4620_ADDRA[5], _7I4614_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_323_4 (_7I4614_$1I4488_$1I4620_ADDRA[4], _7I4614_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_323_3 (_7I4614_$1I4488_$1I4620_ADDRA[3], _7I4614_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_323_2 (_7I4614_$1I4488_$1I4620_ADDRA[2], _7I4614_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_323_1 (_7I4614_$1I4488_$1I4620_ADDRA[1], _7I4614_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_323_0 (_7I4614_$1I4488_$1I4620_ADDRA[0], _7I4614_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _7I4614_$1I4488_$1I4620_ADDRB;
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_324_9 (_7I4614_$1I4488_$1I4620_ADDRB[9], _7I4614_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_324_8 (_7I4614_$1I4488_$1I4620_ADDRB[8], _7I4614_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_324_7 (_7I4614_$1I4488_$1I4620_ADDRB[7], _7I4614_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_324_6 (_7I4614_$1I4488_$1I4620_ADDRB[6], _7I4614_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_324_5 (_7I4614_$1I4488_$1I4620_ADDRB[5], _7I4614_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_324_4 (_7I4614_$1I4488_$1I4620_ADDRB[4], _7I4614_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_324_3 (_7I4614_$1I4488_$1I4620_ADDRB[3], _7I4614_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_324_2 (_7I4614_$1I4488_$1I4620_ADDRB[2], _7I4614_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_324_1 (_7I4614_$1I4488_$1I4620_ADDRB[1], _7I4614_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_324_0 (_7I4614_$1I4488_$1I4620_ADDRB[0], _7I4614_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _7I4614_$1I4488_$1I4620_CLKA;
 reg [1:16] _7I4614_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_325 (_7I4614_$1I4488_$1I4620_CLKA, _7I4614_$1I4488_$1I4620_CLKA__vlIN);

 wire  _7I4614_$1I4488_$1I4620_CLKB;
 reg [1:16] _7I4614_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_326 (_7I4614_$1I4488_$1I4620_CLKB, _7I4614_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _7I4614_$1I4488_$1I4620_DIA;
 reg [1:16] _7I4614_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_327_7 (_7I4614_$1I4488_$1I4620_DIA[7], _7I4614_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_327_6 (_7I4614_$1I4488_$1I4620_DIA[6], _7I4614_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_327_5 (_7I4614_$1I4488_$1I4620_DIA[5], _7I4614_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_327_4 (_7I4614_$1I4488_$1I4620_DIA[4], _7I4614_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_327_3 (_7I4614_$1I4488_$1I4620_DIA[3], _7I4614_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_327_2 (_7I4614_$1I4488_$1I4620_DIA[2], _7I4614_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_327_1 (_7I4614_$1I4488_$1I4620_DIA[1], _7I4614_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_327_0 (_7I4614_$1I4488_$1I4620_DIA[0], _7I4614_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _7I4614_$1I4488_$1I4620_DIB;
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_328_15 (_7I4614_$1I4488_$1I4620_DIB[15], _7I4614_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_328_14 (_7I4614_$1I4488_$1I4620_DIB[14], _7I4614_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_328_13 (_7I4614_$1I4488_$1I4620_DIB[13], _7I4614_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_328_12 (_7I4614_$1I4488_$1I4620_DIB[12], _7I4614_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_328_11 (_7I4614_$1I4488_$1I4620_DIB[11], _7I4614_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_328_10 (_7I4614_$1I4488_$1I4620_DIB[10], _7I4614_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_328_9 (_7I4614_$1I4488_$1I4620_DIB[9], _7I4614_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_328_8 (_7I4614_$1I4488_$1I4620_DIB[8], _7I4614_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_328_7 (_7I4614_$1I4488_$1I4620_DIB[7], _7I4614_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_328_6 (_7I4614_$1I4488_$1I4620_DIB[6], _7I4614_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_328_5 (_7I4614_$1I4488_$1I4620_DIB[5], _7I4614_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_328_4 (_7I4614_$1I4488_$1I4620_DIB[4], _7I4614_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_328_3 (_7I4614_$1I4488_$1I4620_DIB[3], _7I4614_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_328_2 (_7I4614_$1I4488_$1I4620_DIB[2], _7I4614_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_328_1 (_7I4614_$1I4488_$1I4620_DIB[1], _7I4614_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_328_0 (_7I4614_$1I4488_$1I4620_DIB[0], _7I4614_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _7I4614_$1I4488_$1I4620_DIPA;
 reg [1:16] _7I4614_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_329_0 (_7I4614_$1I4488_$1I4620_DIPA[0], _7I4614_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _7I4614_$1I4488_$1I4620_DIPB;
 reg [1:16] _7I4614_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_330_1 (_7I4614_$1I4488_$1I4620_DIPB[1], _7I4614_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _7I4614_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_330_0 (_7I4614_$1I4488_$1I4620_DIPB[0], _7I4614_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _7I4614_$1I4488_$1I4620_ENA;
 reg [1:16] _7I4614_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_331 (_7I4614_$1I4488_$1I4620_ENA, _7I4614_$1I4488_$1I4620_ENA__vlIN);

 wire  _7I4614_$1I4488_$1I4620_ENB;
 reg [1:16] _7I4614_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_332 (_7I4614_$1I4488_$1I4620_ENB, _7I4614_$1I4488_$1I4620_ENB__vlIN);

 wire  _7I4614_$1I4488_$1I4620_SSRA;
 reg [1:16] _7I4614_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_333 (_7I4614_$1I4488_$1I4620_SSRA, _7I4614_$1I4488_$1I4620_SSRA__vlIN);

 wire  _7I4614_$1I4488_$1I4620_SSRB;
 reg [1:16] _7I4614_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_334 (_7I4614_$1I4488_$1I4620_SSRB, _7I4614_$1I4488_$1I4620_SSRB__vlIN);

 wire  _7I4614_$1I4488_$1I4620_WEA;
 reg [1:16] _7I4614_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_335 (_7I4614_$1I4488_$1I4620_WEA, _7I4614_$1I4488_$1I4620_WEA__vlIN);

 wire  _7I4614_$1I4488_$1I4620_WEB;
 reg [1:16] _7I4614_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_336 (_7I4614_$1I4488_$1I4620_WEB, _7I4614_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _7I4614_$1I4488_$1I4620 ( _7I4614_$1I4488_$1I4620_DOA , _7I4614_$1I4488_$1I4620_DOB , _7I4614_$1I4488_$1I4620_DOPA , _7I4614_$1I4488_$1I4620_DOPB , _7I4614_$1I4488_$1I4620_ADDRA , _7I4614_$1I4488_$1I4620_ADDRB , _7I4614_$1I4488_$1I4620_CLKA , _7I4614_$1I4488_$1I4620_CLKB , _7I4614_$1I4488_$1I4620_DIA , _7I4614_$1I4488_$1I4620_DIB , _7I4614_$1I4488_$1I4620_DIPA , _7I4614_$1I4488_$1I4620_DIPB , _7I4614_$1I4488_$1I4620_ENA , _7I4614_$1I4488_$1I4620_ENB , _7I4614_$1I4488_$1I4620_SSRA , _7I4614_$1I4488_$1I4620_SSRB , _7I4614_$1I4488_$1I4620_WEA , _7I4614_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4686_$1I4488_$1I4621_DOA;

 wire [15:0] _6I4686_$1I4488_$1I4621_DOB;

 wire [0:0] _6I4686_$1I4488_$1I4621_DOPA;

 wire [1:0] _6I4686_$1I4488_$1I4621_DOPB;

 wire [10:0] _6I4686_$1I4488_$1I4621_ADDRA;
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_337_10 (_6I4686_$1I4488_$1I4621_ADDRA[10], _6I4686_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_337_9 (_6I4686_$1I4488_$1I4621_ADDRA[9], _6I4686_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_337_8 (_6I4686_$1I4488_$1I4621_ADDRA[8], _6I4686_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_337_7 (_6I4686_$1I4488_$1I4621_ADDRA[7], _6I4686_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_337_6 (_6I4686_$1I4488_$1I4621_ADDRA[6], _6I4686_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_337_5 (_6I4686_$1I4488_$1I4621_ADDRA[5], _6I4686_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_337_4 (_6I4686_$1I4488_$1I4621_ADDRA[4], _6I4686_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_337_3 (_6I4686_$1I4488_$1I4621_ADDRA[3], _6I4686_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_337_2 (_6I4686_$1I4488_$1I4621_ADDRA[2], _6I4686_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_337_1 (_6I4686_$1I4488_$1I4621_ADDRA[1], _6I4686_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_337_0 (_6I4686_$1I4488_$1I4621_ADDRA[0], _6I4686_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _6I4686_$1I4488_$1I4621_ADDRB;
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_338_9 (_6I4686_$1I4488_$1I4621_ADDRB[9], _6I4686_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_338_8 (_6I4686_$1I4488_$1I4621_ADDRB[8], _6I4686_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_338_7 (_6I4686_$1I4488_$1I4621_ADDRB[7], _6I4686_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_338_6 (_6I4686_$1I4488_$1I4621_ADDRB[6], _6I4686_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_338_5 (_6I4686_$1I4488_$1I4621_ADDRB[5], _6I4686_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_338_4 (_6I4686_$1I4488_$1I4621_ADDRB[4], _6I4686_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_338_3 (_6I4686_$1I4488_$1I4621_ADDRB[3], _6I4686_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_338_2 (_6I4686_$1I4488_$1I4621_ADDRB[2], _6I4686_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_338_1 (_6I4686_$1I4488_$1I4621_ADDRB[1], _6I4686_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_338_0 (_6I4686_$1I4488_$1I4621_ADDRB[0], _6I4686_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _6I4686_$1I4488_$1I4621_CLKA;
 reg [1:16] _6I4686_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_339 (_6I4686_$1I4488_$1I4621_CLKA, _6I4686_$1I4488_$1I4621_CLKA__vlIN);

 wire  _6I4686_$1I4488_$1I4621_CLKB;
 reg [1:16] _6I4686_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_340 (_6I4686_$1I4488_$1I4621_CLKB, _6I4686_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _6I4686_$1I4488_$1I4621_DIA;
 reg [1:16] _6I4686_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_341_7 (_6I4686_$1I4488_$1I4621_DIA[7], _6I4686_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_341_6 (_6I4686_$1I4488_$1I4621_DIA[6], _6I4686_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_341_5 (_6I4686_$1I4488_$1I4621_DIA[5], _6I4686_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_341_4 (_6I4686_$1I4488_$1I4621_DIA[4], _6I4686_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_341_3 (_6I4686_$1I4488_$1I4621_DIA[3], _6I4686_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_341_2 (_6I4686_$1I4488_$1I4621_DIA[2], _6I4686_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_341_1 (_6I4686_$1I4488_$1I4621_DIA[1], _6I4686_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_341_0 (_6I4686_$1I4488_$1I4621_DIA[0], _6I4686_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _6I4686_$1I4488_$1I4621_DIB;
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_342_15 (_6I4686_$1I4488_$1I4621_DIB[15], _6I4686_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_342_14 (_6I4686_$1I4488_$1I4621_DIB[14], _6I4686_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_342_13 (_6I4686_$1I4488_$1I4621_DIB[13], _6I4686_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_342_12 (_6I4686_$1I4488_$1I4621_DIB[12], _6I4686_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_342_11 (_6I4686_$1I4488_$1I4621_DIB[11], _6I4686_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_342_10 (_6I4686_$1I4488_$1I4621_DIB[10], _6I4686_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_342_9 (_6I4686_$1I4488_$1I4621_DIB[9], _6I4686_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_342_8 (_6I4686_$1I4488_$1I4621_DIB[8], _6I4686_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_342_7 (_6I4686_$1I4488_$1I4621_DIB[7], _6I4686_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_342_6 (_6I4686_$1I4488_$1I4621_DIB[6], _6I4686_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_342_5 (_6I4686_$1I4488_$1I4621_DIB[5], _6I4686_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_342_4 (_6I4686_$1I4488_$1I4621_DIB[4], _6I4686_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_342_3 (_6I4686_$1I4488_$1I4621_DIB[3], _6I4686_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_342_2 (_6I4686_$1I4488_$1I4621_DIB[2], _6I4686_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_342_1 (_6I4686_$1I4488_$1I4621_DIB[1], _6I4686_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_342_0 (_6I4686_$1I4488_$1I4621_DIB[0], _6I4686_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _6I4686_$1I4488_$1I4621_DIPA;
 reg [1:16] _6I4686_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_343_0 (_6I4686_$1I4488_$1I4621_DIPA[0], _6I4686_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _6I4686_$1I4488_$1I4621_DIPB;
 reg [1:16] _6I4686_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_344_1 (_6I4686_$1I4488_$1I4621_DIPB[1], _6I4686_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_344_0 (_6I4686_$1I4488_$1I4621_DIPB[0], _6I4686_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _6I4686_$1I4488_$1I4621_ENA;
 reg [1:16] _6I4686_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_345 (_6I4686_$1I4488_$1I4621_ENA, _6I4686_$1I4488_$1I4621_ENA__vlIN);

 wire  _6I4686_$1I4488_$1I4621_ENB;
 reg [1:16] _6I4686_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_346 (_6I4686_$1I4488_$1I4621_ENB, _6I4686_$1I4488_$1I4621_ENB__vlIN);

 wire  _6I4686_$1I4488_$1I4621_SSRA;
 reg [1:16] _6I4686_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_347 (_6I4686_$1I4488_$1I4621_SSRA, _6I4686_$1I4488_$1I4621_SSRA__vlIN);

 wire  _6I4686_$1I4488_$1I4621_SSRB;
 reg [1:16] _6I4686_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_348 (_6I4686_$1I4488_$1I4621_SSRB, _6I4686_$1I4488_$1I4621_SSRB__vlIN);

 wire  _6I4686_$1I4488_$1I4621_WEA;
 reg [1:16] _6I4686_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_349 (_6I4686_$1I4488_$1I4621_WEA, _6I4686_$1I4488_$1I4621_WEA__vlIN);

 wire  _6I4686_$1I4488_$1I4621_WEB;
 reg [1:16] _6I4686_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_350 (_6I4686_$1I4488_$1I4621_WEB, _6I4686_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _6I4686_$1I4488_$1I4621 ( _6I4686_$1I4488_$1I4621_DOA , _6I4686_$1I4488_$1I4621_DOB , _6I4686_$1I4488_$1I4621_DOPA , _6I4686_$1I4488_$1I4621_DOPB , _6I4686_$1I4488_$1I4621_ADDRA , _6I4686_$1I4488_$1I4621_ADDRB , _6I4686_$1I4488_$1I4621_CLKA , _6I4686_$1I4488_$1I4621_CLKB , _6I4686_$1I4488_$1I4621_DIA , _6I4686_$1I4488_$1I4621_DIB , _6I4686_$1I4488_$1I4621_DIPA , _6I4686_$1I4488_$1I4621_DIPB , _6I4686_$1I4488_$1I4621_ENA , _6I4686_$1I4488_$1I4621_ENB , _6I4686_$1I4488_$1I4621_SSRA , _6I4686_$1I4488_$1I4621_SSRB , _6I4686_$1I4488_$1I4621_WEA , _6I4686_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4686_$1I4488_$1I4620_DOA;

 wire [15:0] _6I4686_$1I4488_$1I4620_DOB;

 wire [0:0] _6I4686_$1I4488_$1I4620_DOPA;

 wire [1:0] _6I4686_$1I4488_$1I4620_DOPB;

 wire [10:0] _6I4686_$1I4488_$1I4620_ADDRA;
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_351_10 (_6I4686_$1I4488_$1I4620_ADDRA[10], _6I4686_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_351_9 (_6I4686_$1I4488_$1I4620_ADDRA[9], _6I4686_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_351_8 (_6I4686_$1I4488_$1I4620_ADDRA[8], _6I4686_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_351_7 (_6I4686_$1I4488_$1I4620_ADDRA[7], _6I4686_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_351_6 (_6I4686_$1I4488_$1I4620_ADDRA[6], _6I4686_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_351_5 (_6I4686_$1I4488_$1I4620_ADDRA[5], _6I4686_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_351_4 (_6I4686_$1I4488_$1I4620_ADDRA[4], _6I4686_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_351_3 (_6I4686_$1I4488_$1I4620_ADDRA[3], _6I4686_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_351_2 (_6I4686_$1I4488_$1I4620_ADDRA[2], _6I4686_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_351_1 (_6I4686_$1I4488_$1I4620_ADDRA[1], _6I4686_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_351_0 (_6I4686_$1I4488_$1I4620_ADDRA[0], _6I4686_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _6I4686_$1I4488_$1I4620_ADDRB;
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_352_9 (_6I4686_$1I4488_$1I4620_ADDRB[9], _6I4686_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_352_8 (_6I4686_$1I4488_$1I4620_ADDRB[8], _6I4686_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_352_7 (_6I4686_$1I4488_$1I4620_ADDRB[7], _6I4686_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_352_6 (_6I4686_$1I4488_$1I4620_ADDRB[6], _6I4686_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_352_5 (_6I4686_$1I4488_$1I4620_ADDRB[5], _6I4686_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_352_4 (_6I4686_$1I4488_$1I4620_ADDRB[4], _6I4686_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_352_3 (_6I4686_$1I4488_$1I4620_ADDRB[3], _6I4686_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_352_2 (_6I4686_$1I4488_$1I4620_ADDRB[2], _6I4686_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_352_1 (_6I4686_$1I4488_$1I4620_ADDRB[1], _6I4686_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_352_0 (_6I4686_$1I4488_$1I4620_ADDRB[0], _6I4686_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _6I4686_$1I4488_$1I4620_CLKA;
 reg [1:16] _6I4686_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_353 (_6I4686_$1I4488_$1I4620_CLKA, _6I4686_$1I4488_$1I4620_CLKA__vlIN);

 wire  _6I4686_$1I4488_$1I4620_CLKB;
 reg [1:16] _6I4686_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_354 (_6I4686_$1I4488_$1I4620_CLKB, _6I4686_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _6I4686_$1I4488_$1I4620_DIA;
 reg [1:16] _6I4686_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_355_7 (_6I4686_$1I4488_$1I4620_DIA[7], _6I4686_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_355_6 (_6I4686_$1I4488_$1I4620_DIA[6], _6I4686_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_355_5 (_6I4686_$1I4488_$1I4620_DIA[5], _6I4686_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_355_4 (_6I4686_$1I4488_$1I4620_DIA[4], _6I4686_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_355_3 (_6I4686_$1I4488_$1I4620_DIA[3], _6I4686_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_355_2 (_6I4686_$1I4488_$1I4620_DIA[2], _6I4686_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_355_1 (_6I4686_$1I4488_$1I4620_DIA[1], _6I4686_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_355_0 (_6I4686_$1I4488_$1I4620_DIA[0], _6I4686_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _6I4686_$1I4488_$1I4620_DIB;
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_356_15 (_6I4686_$1I4488_$1I4620_DIB[15], _6I4686_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_356_14 (_6I4686_$1I4488_$1I4620_DIB[14], _6I4686_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_356_13 (_6I4686_$1I4488_$1I4620_DIB[13], _6I4686_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_356_12 (_6I4686_$1I4488_$1I4620_DIB[12], _6I4686_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_356_11 (_6I4686_$1I4488_$1I4620_DIB[11], _6I4686_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_356_10 (_6I4686_$1I4488_$1I4620_DIB[10], _6I4686_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_356_9 (_6I4686_$1I4488_$1I4620_DIB[9], _6I4686_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_356_8 (_6I4686_$1I4488_$1I4620_DIB[8], _6I4686_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_356_7 (_6I4686_$1I4488_$1I4620_DIB[7], _6I4686_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_356_6 (_6I4686_$1I4488_$1I4620_DIB[6], _6I4686_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_356_5 (_6I4686_$1I4488_$1I4620_DIB[5], _6I4686_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_356_4 (_6I4686_$1I4488_$1I4620_DIB[4], _6I4686_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_356_3 (_6I4686_$1I4488_$1I4620_DIB[3], _6I4686_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_356_2 (_6I4686_$1I4488_$1I4620_DIB[2], _6I4686_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_356_1 (_6I4686_$1I4488_$1I4620_DIB[1], _6I4686_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_356_0 (_6I4686_$1I4488_$1I4620_DIB[0], _6I4686_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _6I4686_$1I4488_$1I4620_DIPA;
 reg [1:16] _6I4686_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_357_0 (_6I4686_$1I4488_$1I4620_DIPA[0], _6I4686_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _6I4686_$1I4488_$1I4620_DIPB;
 reg [1:16] _6I4686_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_358_1 (_6I4686_$1I4488_$1I4620_DIPB[1], _6I4686_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _6I4686_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_358_0 (_6I4686_$1I4488_$1I4620_DIPB[0], _6I4686_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _6I4686_$1I4488_$1I4620_ENA;
 reg [1:16] _6I4686_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_359 (_6I4686_$1I4488_$1I4620_ENA, _6I4686_$1I4488_$1I4620_ENA__vlIN);

 wire  _6I4686_$1I4488_$1I4620_ENB;
 reg [1:16] _6I4686_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_360 (_6I4686_$1I4488_$1I4620_ENB, _6I4686_$1I4488_$1I4620_ENB__vlIN);

 wire  _6I4686_$1I4488_$1I4620_SSRA;
 reg [1:16] _6I4686_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_361 (_6I4686_$1I4488_$1I4620_SSRA, _6I4686_$1I4488_$1I4620_SSRA__vlIN);

 wire  _6I4686_$1I4488_$1I4620_SSRB;
 reg [1:16] _6I4686_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_362 (_6I4686_$1I4488_$1I4620_SSRB, _6I4686_$1I4488_$1I4620_SSRB__vlIN);

 wire  _6I4686_$1I4488_$1I4620_WEA;
 reg [1:16] _6I4686_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_363 (_6I4686_$1I4488_$1I4620_WEA, _6I4686_$1I4488_$1I4620_WEA__vlIN);

 wire  _6I4686_$1I4488_$1I4620_WEB;
 reg [1:16] _6I4686_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_364 (_6I4686_$1I4488_$1I4620_WEB, _6I4686_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _6I4686_$1I4488_$1I4620 ( _6I4686_$1I4488_$1I4620_DOA , _6I4686_$1I4488_$1I4620_DOB , _6I4686_$1I4488_$1I4620_DOPA , _6I4686_$1I4488_$1I4620_DOPB , _6I4686_$1I4488_$1I4620_ADDRA , _6I4686_$1I4488_$1I4620_ADDRB , _6I4686_$1I4488_$1I4620_CLKA , _6I4686_$1I4488_$1I4620_CLKB , _6I4686_$1I4488_$1I4620_DIA , _6I4686_$1I4488_$1I4620_DIB , _6I4686_$1I4488_$1I4620_DIPA , _6I4686_$1I4488_$1I4620_DIPB , _6I4686_$1I4488_$1I4620_ENA , _6I4686_$1I4488_$1I4620_ENB , _6I4686_$1I4488_$1I4620_SSRA , _6I4686_$1I4488_$1I4620_SSRB , _6I4686_$1I4488_$1I4620_WEA , _6I4686_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4641_$1I4488_$1I4621_DOA;

 wire [15:0] _6I4641_$1I4488_$1I4621_DOB;

 wire [0:0] _6I4641_$1I4488_$1I4621_DOPA;

 wire [1:0] _6I4641_$1I4488_$1I4621_DOPB;

 wire [10:0] _6I4641_$1I4488_$1I4621_ADDRA;
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_365_10 (_6I4641_$1I4488_$1I4621_ADDRA[10], _6I4641_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_365_9 (_6I4641_$1I4488_$1I4621_ADDRA[9], _6I4641_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_365_8 (_6I4641_$1I4488_$1I4621_ADDRA[8], _6I4641_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_365_7 (_6I4641_$1I4488_$1I4621_ADDRA[7], _6I4641_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_365_6 (_6I4641_$1I4488_$1I4621_ADDRA[6], _6I4641_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_365_5 (_6I4641_$1I4488_$1I4621_ADDRA[5], _6I4641_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_365_4 (_6I4641_$1I4488_$1I4621_ADDRA[4], _6I4641_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_365_3 (_6I4641_$1I4488_$1I4621_ADDRA[3], _6I4641_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_365_2 (_6I4641_$1I4488_$1I4621_ADDRA[2], _6I4641_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_365_1 (_6I4641_$1I4488_$1I4621_ADDRA[1], _6I4641_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_365_0 (_6I4641_$1I4488_$1I4621_ADDRA[0], _6I4641_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _6I4641_$1I4488_$1I4621_ADDRB;
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_366_9 (_6I4641_$1I4488_$1I4621_ADDRB[9], _6I4641_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_366_8 (_6I4641_$1I4488_$1I4621_ADDRB[8], _6I4641_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_366_7 (_6I4641_$1I4488_$1I4621_ADDRB[7], _6I4641_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_366_6 (_6I4641_$1I4488_$1I4621_ADDRB[6], _6I4641_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_366_5 (_6I4641_$1I4488_$1I4621_ADDRB[5], _6I4641_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_366_4 (_6I4641_$1I4488_$1I4621_ADDRB[4], _6I4641_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_366_3 (_6I4641_$1I4488_$1I4621_ADDRB[3], _6I4641_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_366_2 (_6I4641_$1I4488_$1I4621_ADDRB[2], _6I4641_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_366_1 (_6I4641_$1I4488_$1I4621_ADDRB[1], _6I4641_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_366_0 (_6I4641_$1I4488_$1I4621_ADDRB[0], _6I4641_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _6I4641_$1I4488_$1I4621_CLKA;
 reg [1:16] _6I4641_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_367 (_6I4641_$1I4488_$1I4621_CLKA, _6I4641_$1I4488_$1I4621_CLKA__vlIN);

 wire  _6I4641_$1I4488_$1I4621_CLKB;
 reg [1:16] _6I4641_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_368 (_6I4641_$1I4488_$1I4621_CLKB, _6I4641_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _6I4641_$1I4488_$1I4621_DIA;
 reg [1:16] _6I4641_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_369_7 (_6I4641_$1I4488_$1I4621_DIA[7], _6I4641_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_369_6 (_6I4641_$1I4488_$1I4621_DIA[6], _6I4641_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_369_5 (_6I4641_$1I4488_$1I4621_DIA[5], _6I4641_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_369_4 (_6I4641_$1I4488_$1I4621_DIA[4], _6I4641_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_369_3 (_6I4641_$1I4488_$1I4621_DIA[3], _6I4641_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_369_2 (_6I4641_$1I4488_$1I4621_DIA[2], _6I4641_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_369_1 (_6I4641_$1I4488_$1I4621_DIA[1], _6I4641_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_369_0 (_6I4641_$1I4488_$1I4621_DIA[0], _6I4641_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _6I4641_$1I4488_$1I4621_DIB;
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_370_15 (_6I4641_$1I4488_$1I4621_DIB[15], _6I4641_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_370_14 (_6I4641_$1I4488_$1I4621_DIB[14], _6I4641_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_370_13 (_6I4641_$1I4488_$1I4621_DIB[13], _6I4641_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_370_12 (_6I4641_$1I4488_$1I4621_DIB[12], _6I4641_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_370_11 (_6I4641_$1I4488_$1I4621_DIB[11], _6I4641_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_370_10 (_6I4641_$1I4488_$1I4621_DIB[10], _6I4641_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_370_9 (_6I4641_$1I4488_$1I4621_DIB[9], _6I4641_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_370_8 (_6I4641_$1I4488_$1I4621_DIB[8], _6I4641_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_370_7 (_6I4641_$1I4488_$1I4621_DIB[7], _6I4641_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_370_6 (_6I4641_$1I4488_$1I4621_DIB[6], _6I4641_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_370_5 (_6I4641_$1I4488_$1I4621_DIB[5], _6I4641_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_370_4 (_6I4641_$1I4488_$1I4621_DIB[4], _6I4641_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_370_3 (_6I4641_$1I4488_$1I4621_DIB[3], _6I4641_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_370_2 (_6I4641_$1I4488_$1I4621_DIB[2], _6I4641_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_370_1 (_6I4641_$1I4488_$1I4621_DIB[1], _6I4641_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_370_0 (_6I4641_$1I4488_$1I4621_DIB[0], _6I4641_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _6I4641_$1I4488_$1I4621_DIPA;
 reg [1:16] _6I4641_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_371_0 (_6I4641_$1I4488_$1I4621_DIPA[0], _6I4641_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _6I4641_$1I4488_$1I4621_DIPB;
 reg [1:16] _6I4641_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_372_1 (_6I4641_$1I4488_$1I4621_DIPB[1], _6I4641_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_372_0 (_6I4641_$1I4488_$1I4621_DIPB[0], _6I4641_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _6I4641_$1I4488_$1I4621_ENA;
 reg [1:16] _6I4641_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_373 (_6I4641_$1I4488_$1I4621_ENA, _6I4641_$1I4488_$1I4621_ENA__vlIN);

 wire  _6I4641_$1I4488_$1I4621_ENB;
 reg [1:16] _6I4641_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_374 (_6I4641_$1I4488_$1I4621_ENB, _6I4641_$1I4488_$1I4621_ENB__vlIN);

 wire  _6I4641_$1I4488_$1I4621_SSRA;
 reg [1:16] _6I4641_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_375 (_6I4641_$1I4488_$1I4621_SSRA, _6I4641_$1I4488_$1I4621_SSRA__vlIN);

 wire  _6I4641_$1I4488_$1I4621_SSRB;
 reg [1:16] _6I4641_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_376 (_6I4641_$1I4488_$1I4621_SSRB, _6I4641_$1I4488_$1I4621_SSRB__vlIN);

 wire  _6I4641_$1I4488_$1I4621_WEA;
 reg [1:16] _6I4641_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_377 (_6I4641_$1I4488_$1I4621_WEA, _6I4641_$1I4488_$1I4621_WEA__vlIN);

 wire  _6I4641_$1I4488_$1I4621_WEB;
 reg [1:16] _6I4641_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_378 (_6I4641_$1I4488_$1I4621_WEB, _6I4641_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _6I4641_$1I4488_$1I4621 ( _6I4641_$1I4488_$1I4621_DOA , _6I4641_$1I4488_$1I4621_DOB , _6I4641_$1I4488_$1I4621_DOPA , _6I4641_$1I4488_$1I4621_DOPB , _6I4641_$1I4488_$1I4621_ADDRA , _6I4641_$1I4488_$1I4621_ADDRB , _6I4641_$1I4488_$1I4621_CLKA , _6I4641_$1I4488_$1I4621_CLKB , _6I4641_$1I4488_$1I4621_DIA , _6I4641_$1I4488_$1I4621_DIB , _6I4641_$1I4488_$1I4621_DIPA , _6I4641_$1I4488_$1I4621_DIPB , _6I4641_$1I4488_$1I4621_ENA , _6I4641_$1I4488_$1I4621_ENB , _6I4641_$1I4488_$1I4621_SSRA , _6I4641_$1I4488_$1I4621_SSRB , _6I4641_$1I4488_$1I4621_WEA , _6I4641_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4641_$1I4488_$1I4620_DOA;

 wire [15:0] _6I4641_$1I4488_$1I4620_DOB;

 wire [0:0] _6I4641_$1I4488_$1I4620_DOPA;

 wire [1:0] _6I4641_$1I4488_$1I4620_DOPB;

 wire [10:0] _6I4641_$1I4488_$1I4620_ADDRA;
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_379_10 (_6I4641_$1I4488_$1I4620_ADDRA[10], _6I4641_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_379_9 (_6I4641_$1I4488_$1I4620_ADDRA[9], _6I4641_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_379_8 (_6I4641_$1I4488_$1I4620_ADDRA[8], _6I4641_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_379_7 (_6I4641_$1I4488_$1I4620_ADDRA[7], _6I4641_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_379_6 (_6I4641_$1I4488_$1I4620_ADDRA[6], _6I4641_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_379_5 (_6I4641_$1I4488_$1I4620_ADDRA[5], _6I4641_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_379_4 (_6I4641_$1I4488_$1I4620_ADDRA[4], _6I4641_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_379_3 (_6I4641_$1I4488_$1I4620_ADDRA[3], _6I4641_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_379_2 (_6I4641_$1I4488_$1I4620_ADDRA[2], _6I4641_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_379_1 (_6I4641_$1I4488_$1I4620_ADDRA[1], _6I4641_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_379_0 (_6I4641_$1I4488_$1I4620_ADDRA[0], _6I4641_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _6I4641_$1I4488_$1I4620_ADDRB;
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_380_9 (_6I4641_$1I4488_$1I4620_ADDRB[9], _6I4641_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_380_8 (_6I4641_$1I4488_$1I4620_ADDRB[8], _6I4641_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_380_7 (_6I4641_$1I4488_$1I4620_ADDRB[7], _6I4641_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_380_6 (_6I4641_$1I4488_$1I4620_ADDRB[6], _6I4641_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_380_5 (_6I4641_$1I4488_$1I4620_ADDRB[5], _6I4641_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_380_4 (_6I4641_$1I4488_$1I4620_ADDRB[4], _6I4641_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_380_3 (_6I4641_$1I4488_$1I4620_ADDRB[3], _6I4641_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_380_2 (_6I4641_$1I4488_$1I4620_ADDRB[2], _6I4641_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_380_1 (_6I4641_$1I4488_$1I4620_ADDRB[1], _6I4641_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_380_0 (_6I4641_$1I4488_$1I4620_ADDRB[0], _6I4641_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _6I4641_$1I4488_$1I4620_CLKA;
 reg [1:16] _6I4641_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_381 (_6I4641_$1I4488_$1I4620_CLKA, _6I4641_$1I4488_$1I4620_CLKA__vlIN);

 wire  _6I4641_$1I4488_$1I4620_CLKB;
 reg [1:16] _6I4641_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_382 (_6I4641_$1I4488_$1I4620_CLKB, _6I4641_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _6I4641_$1I4488_$1I4620_DIA;
 reg [1:16] _6I4641_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_383_7 (_6I4641_$1I4488_$1I4620_DIA[7], _6I4641_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_383_6 (_6I4641_$1I4488_$1I4620_DIA[6], _6I4641_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_383_5 (_6I4641_$1I4488_$1I4620_DIA[5], _6I4641_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_383_4 (_6I4641_$1I4488_$1I4620_DIA[4], _6I4641_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_383_3 (_6I4641_$1I4488_$1I4620_DIA[3], _6I4641_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_383_2 (_6I4641_$1I4488_$1I4620_DIA[2], _6I4641_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_383_1 (_6I4641_$1I4488_$1I4620_DIA[1], _6I4641_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_383_0 (_6I4641_$1I4488_$1I4620_DIA[0], _6I4641_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _6I4641_$1I4488_$1I4620_DIB;
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_384_15 (_6I4641_$1I4488_$1I4620_DIB[15], _6I4641_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_384_14 (_6I4641_$1I4488_$1I4620_DIB[14], _6I4641_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_384_13 (_6I4641_$1I4488_$1I4620_DIB[13], _6I4641_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_384_12 (_6I4641_$1I4488_$1I4620_DIB[12], _6I4641_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_384_11 (_6I4641_$1I4488_$1I4620_DIB[11], _6I4641_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_384_10 (_6I4641_$1I4488_$1I4620_DIB[10], _6I4641_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_384_9 (_6I4641_$1I4488_$1I4620_DIB[9], _6I4641_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_384_8 (_6I4641_$1I4488_$1I4620_DIB[8], _6I4641_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_384_7 (_6I4641_$1I4488_$1I4620_DIB[7], _6I4641_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_384_6 (_6I4641_$1I4488_$1I4620_DIB[6], _6I4641_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_384_5 (_6I4641_$1I4488_$1I4620_DIB[5], _6I4641_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_384_4 (_6I4641_$1I4488_$1I4620_DIB[4], _6I4641_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_384_3 (_6I4641_$1I4488_$1I4620_DIB[3], _6I4641_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_384_2 (_6I4641_$1I4488_$1I4620_DIB[2], _6I4641_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_384_1 (_6I4641_$1I4488_$1I4620_DIB[1], _6I4641_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_384_0 (_6I4641_$1I4488_$1I4620_DIB[0], _6I4641_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _6I4641_$1I4488_$1I4620_DIPA;
 reg [1:16] _6I4641_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_385_0 (_6I4641_$1I4488_$1I4620_DIPA[0], _6I4641_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _6I4641_$1I4488_$1I4620_DIPB;
 reg [1:16] _6I4641_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_386_1 (_6I4641_$1I4488_$1I4620_DIPB[1], _6I4641_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _6I4641_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_386_0 (_6I4641_$1I4488_$1I4620_DIPB[0], _6I4641_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _6I4641_$1I4488_$1I4620_ENA;
 reg [1:16] _6I4641_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_387 (_6I4641_$1I4488_$1I4620_ENA, _6I4641_$1I4488_$1I4620_ENA__vlIN);

 wire  _6I4641_$1I4488_$1I4620_ENB;
 reg [1:16] _6I4641_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_388 (_6I4641_$1I4488_$1I4620_ENB, _6I4641_$1I4488_$1I4620_ENB__vlIN);

 wire  _6I4641_$1I4488_$1I4620_SSRA;
 reg [1:16] _6I4641_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_389 (_6I4641_$1I4488_$1I4620_SSRA, _6I4641_$1I4488_$1I4620_SSRA__vlIN);

 wire  _6I4641_$1I4488_$1I4620_SSRB;
 reg [1:16] _6I4641_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_390 (_6I4641_$1I4488_$1I4620_SSRB, _6I4641_$1I4488_$1I4620_SSRB__vlIN);

 wire  _6I4641_$1I4488_$1I4620_WEA;
 reg [1:16] _6I4641_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_391 (_6I4641_$1I4488_$1I4620_WEA, _6I4641_$1I4488_$1I4620_WEA__vlIN);

 wire  _6I4641_$1I4488_$1I4620_WEB;
 reg [1:16] _6I4641_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_392 (_6I4641_$1I4488_$1I4620_WEB, _6I4641_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _6I4641_$1I4488_$1I4620 ( _6I4641_$1I4488_$1I4620_DOA , _6I4641_$1I4488_$1I4620_DOB , _6I4641_$1I4488_$1I4620_DOPA , _6I4641_$1I4488_$1I4620_DOPB , _6I4641_$1I4488_$1I4620_ADDRA , _6I4641_$1I4488_$1I4620_ADDRB , _6I4641_$1I4488_$1I4620_CLKA , _6I4641_$1I4488_$1I4620_CLKB , _6I4641_$1I4488_$1I4620_DIA , _6I4641_$1I4488_$1I4620_DIB , _6I4641_$1I4488_$1I4620_DIPA , _6I4641_$1I4488_$1I4620_DIPB , _6I4641_$1I4488_$1I4620_ENA , _6I4641_$1I4488_$1I4620_ENB , _6I4641_$1I4488_$1I4620_SSRA , _6I4641_$1I4488_$1I4620_SSRB , _6I4641_$1I4488_$1I4620_WEA , _6I4641_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4614_$1I4488_$1I4621_DOA;

 wire [15:0] _6I4614_$1I4488_$1I4621_DOB;

 wire [0:0] _6I4614_$1I4488_$1I4621_DOPA;

 wire [1:0] _6I4614_$1I4488_$1I4621_DOPB;

 wire [10:0] _6I4614_$1I4488_$1I4621_ADDRA;
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_393_10 (_6I4614_$1I4488_$1I4621_ADDRA[10], _6I4614_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_393_9 (_6I4614_$1I4488_$1I4621_ADDRA[9], _6I4614_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_393_8 (_6I4614_$1I4488_$1I4621_ADDRA[8], _6I4614_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_393_7 (_6I4614_$1I4488_$1I4621_ADDRA[7], _6I4614_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_393_6 (_6I4614_$1I4488_$1I4621_ADDRA[6], _6I4614_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_393_5 (_6I4614_$1I4488_$1I4621_ADDRA[5], _6I4614_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_393_4 (_6I4614_$1I4488_$1I4621_ADDRA[4], _6I4614_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_393_3 (_6I4614_$1I4488_$1I4621_ADDRA[3], _6I4614_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_393_2 (_6I4614_$1I4488_$1I4621_ADDRA[2], _6I4614_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_393_1 (_6I4614_$1I4488_$1I4621_ADDRA[1], _6I4614_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_393_0 (_6I4614_$1I4488_$1I4621_ADDRA[0], _6I4614_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _6I4614_$1I4488_$1I4621_ADDRB;
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_394_9 (_6I4614_$1I4488_$1I4621_ADDRB[9], _6I4614_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_394_8 (_6I4614_$1I4488_$1I4621_ADDRB[8], _6I4614_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_394_7 (_6I4614_$1I4488_$1I4621_ADDRB[7], _6I4614_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_394_6 (_6I4614_$1I4488_$1I4621_ADDRB[6], _6I4614_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_394_5 (_6I4614_$1I4488_$1I4621_ADDRB[5], _6I4614_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_394_4 (_6I4614_$1I4488_$1I4621_ADDRB[4], _6I4614_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_394_3 (_6I4614_$1I4488_$1I4621_ADDRB[3], _6I4614_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_394_2 (_6I4614_$1I4488_$1I4621_ADDRB[2], _6I4614_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_394_1 (_6I4614_$1I4488_$1I4621_ADDRB[1], _6I4614_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_394_0 (_6I4614_$1I4488_$1I4621_ADDRB[0], _6I4614_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _6I4614_$1I4488_$1I4621_CLKA;
 reg [1:16] _6I4614_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_395 (_6I4614_$1I4488_$1I4621_CLKA, _6I4614_$1I4488_$1I4621_CLKA__vlIN);

 wire  _6I4614_$1I4488_$1I4621_CLKB;
 reg [1:16] _6I4614_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_396 (_6I4614_$1I4488_$1I4621_CLKB, _6I4614_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _6I4614_$1I4488_$1I4621_DIA;
 reg [1:16] _6I4614_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_397_7 (_6I4614_$1I4488_$1I4621_DIA[7], _6I4614_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_397_6 (_6I4614_$1I4488_$1I4621_DIA[6], _6I4614_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_397_5 (_6I4614_$1I4488_$1I4621_DIA[5], _6I4614_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_397_4 (_6I4614_$1I4488_$1I4621_DIA[4], _6I4614_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_397_3 (_6I4614_$1I4488_$1I4621_DIA[3], _6I4614_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_397_2 (_6I4614_$1I4488_$1I4621_DIA[2], _6I4614_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_397_1 (_6I4614_$1I4488_$1I4621_DIA[1], _6I4614_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_397_0 (_6I4614_$1I4488_$1I4621_DIA[0], _6I4614_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _6I4614_$1I4488_$1I4621_DIB;
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_398_15 (_6I4614_$1I4488_$1I4621_DIB[15], _6I4614_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_398_14 (_6I4614_$1I4488_$1I4621_DIB[14], _6I4614_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_398_13 (_6I4614_$1I4488_$1I4621_DIB[13], _6I4614_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_398_12 (_6I4614_$1I4488_$1I4621_DIB[12], _6I4614_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_398_11 (_6I4614_$1I4488_$1I4621_DIB[11], _6I4614_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_398_10 (_6I4614_$1I4488_$1I4621_DIB[10], _6I4614_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_398_9 (_6I4614_$1I4488_$1I4621_DIB[9], _6I4614_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_398_8 (_6I4614_$1I4488_$1I4621_DIB[8], _6I4614_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_398_7 (_6I4614_$1I4488_$1I4621_DIB[7], _6I4614_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_398_6 (_6I4614_$1I4488_$1I4621_DIB[6], _6I4614_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_398_5 (_6I4614_$1I4488_$1I4621_DIB[5], _6I4614_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_398_4 (_6I4614_$1I4488_$1I4621_DIB[4], _6I4614_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_398_3 (_6I4614_$1I4488_$1I4621_DIB[3], _6I4614_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_398_2 (_6I4614_$1I4488_$1I4621_DIB[2], _6I4614_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_398_1 (_6I4614_$1I4488_$1I4621_DIB[1], _6I4614_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_398_0 (_6I4614_$1I4488_$1I4621_DIB[0], _6I4614_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _6I4614_$1I4488_$1I4621_DIPA;
 reg [1:16] _6I4614_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_399_0 (_6I4614_$1I4488_$1I4621_DIPA[0], _6I4614_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _6I4614_$1I4488_$1I4621_DIPB;
 reg [1:16] _6I4614_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_400_1 (_6I4614_$1I4488_$1I4621_DIPB[1], _6I4614_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_400_0 (_6I4614_$1I4488_$1I4621_DIPB[0], _6I4614_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _6I4614_$1I4488_$1I4621_ENA;
 reg [1:16] _6I4614_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_401 (_6I4614_$1I4488_$1I4621_ENA, _6I4614_$1I4488_$1I4621_ENA__vlIN);

 wire  _6I4614_$1I4488_$1I4621_ENB;
 reg [1:16] _6I4614_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_402 (_6I4614_$1I4488_$1I4621_ENB, _6I4614_$1I4488_$1I4621_ENB__vlIN);

 wire  _6I4614_$1I4488_$1I4621_SSRA;
 reg [1:16] _6I4614_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_403 (_6I4614_$1I4488_$1I4621_SSRA, _6I4614_$1I4488_$1I4621_SSRA__vlIN);

 wire  _6I4614_$1I4488_$1I4621_SSRB;
 reg [1:16] _6I4614_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_404 (_6I4614_$1I4488_$1I4621_SSRB, _6I4614_$1I4488_$1I4621_SSRB__vlIN);

 wire  _6I4614_$1I4488_$1I4621_WEA;
 reg [1:16] _6I4614_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_405 (_6I4614_$1I4488_$1I4621_WEA, _6I4614_$1I4488_$1I4621_WEA__vlIN);

 wire  _6I4614_$1I4488_$1I4621_WEB;
 reg [1:16] _6I4614_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_406 (_6I4614_$1I4488_$1I4621_WEB, _6I4614_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _6I4614_$1I4488_$1I4621 ( _6I4614_$1I4488_$1I4621_DOA , _6I4614_$1I4488_$1I4621_DOB , _6I4614_$1I4488_$1I4621_DOPA , _6I4614_$1I4488_$1I4621_DOPB , _6I4614_$1I4488_$1I4621_ADDRA , _6I4614_$1I4488_$1I4621_ADDRB , _6I4614_$1I4488_$1I4621_CLKA , _6I4614_$1I4488_$1I4621_CLKB , _6I4614_$1I4488_$1I4621_DIA , _6I4614_$1I4488_$1I4621_DIB , _6I4614_$1I4488_$1I4621_DIPA , _6I4614_$1I4488_$1I4621_DIPB , _6I4614_$1I4488_$1I4621_ENA , _6I4614_$1I4488_$1I4621_ENB , _6I4614_$1I4488_$1I4621_SSRA , _6I4614_$1I4488_$1I4621_SSRB , _6I4614_$1I4488_$1I4621_WEA , _6I4614_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4614_$1I4488_$1I4620_DOA;

 wire [15:0] _6I4614_$1I4488_$1I4620_DOB;

 wire [0:0] _6I4614_$1I4488_$1I4620_DOPA;

 wire [1:0] _6I4614_$1I4488_$1I4620_DOPB;

 wire [10:0] _6I4614_$1I4488_$1I4620_ADDRA;
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_407_10 (_6I4614_$1I4488_$1I4620_ADDRA[10], _6I4614_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_407_9 (_6I4614_$1I4488_$1I4620_ADDRA[9], _6I4614_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_407_8 (_6I4614_$1I4488_$1I4620_ADDRA[8], _6I4614_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_407_7 (_6I4614_$1I4488_$1I4620_ADDRA[7], _6I4614_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_407_6 (_6I4614_$1I4488_$1I4620_ADDRA[6], _6I4614_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_407_5 (_6I4614_$1I4488_$1I4620_ADDRA[5], _6I4614_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_407_4 (_6I4614_$1I4488_$1I4620_ADDRA[4], _6I4614_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_407_3 (_6I4614_$1I4488_$1I4620_ADDRA[3], _6I4614_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_407_2 (_6I4614_$1I4488_$1I4620_ADDRA[2], _6I4614_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_407_1 (_6I4614_$1I4488_$1I4620_ADDRA[1], _6I4614_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_407_0 (_6I4614_$1I4488_$1I4620_ADDRA[0], _6I4614_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _6I4614_$1I4488_$1I4620_ADDRB;
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_408_9 (_6I4614_$1I4488_$1I4620_ADDRB[9], _6I4614_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_408_8 (_6I4614_$1I4488_$1I4620_ADDRB[8], _6I4614_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_408_7 (_6I4614_$1I4488_$1I4620_ADDRB[7], _6I4614_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_408_6 (_6I4614_$1I4488_$1I4620_ADDRB[6], _6I4614_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_408_5 (_6I4614_$1I4488_$1I4620_ADDRB[5], _6I4614_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_408_4 (_6I4614_$1I4488_$1I4620_ADDRB[4], _6I4614_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_408_3 (_6I4614_$1I4488_$1I4620_ADDRB[3], _6I4614_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_408_2 (_6I4614_$1I4488_$1I4620_ADDRB[2], _6I4614_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_408_1 (_6I4614_$1I4488_$1I4620_ADDRB[1], _6I4614_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_408_0 (_6I4614_$1I4488_$1I4620_ADDRB[0], _6I4614_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _6I4614_$1I4488_$1I4620_CLKA;
 reg [1:16] _6I4614_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_409 (_6I4614_$1I4488_$1I4620_CLKA, _6I4614_$1I4488_$1I4620_CLKA__vlIN);

 wire  _6I4614_$1I4488_$1I4620_CLKB;
 reg [1:16] _6I4614_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_410 (_6I4614_$1I4488_$1I4620_CLKB, _6I4614_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _6I4614_$1I4488_$1I4620_DIA;
 reg [1:16] _6I4614_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_411_7 (_6I4614_$1I4488_$1I4620_DIA[7], _6I4614_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_411_6 (_6I4614_$1I4488_$1I4620_DIA[6], _6I4614_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_411_5 (_6I4614_$1I4488_$1I4620_DIA[5], _6I4614_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_411_4 (_6I4614_$1I4488_$1I4620_DIA[4], _6I4614_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_411_3 (_6I4614_$1I4488_$1I4620_DIA[3], _6I4614_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_411_2 (_6I4614_$1I4488_$1I4620_DIA[2], _6I4614_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_411_1 (_6I4614_$1I4488_$1I4620_DIA[1], _6I4614_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_411_0 (_6I4614_$1I4488_$1I4620_DIA[0], _6I4614_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _6I4614_$1I4488_$1I4620_DIB;
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_412_15 (_6I4614_$1I4488_$1I4620_DIB[15], _6I4614_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_412_14 (_6I4614_$1I4488_$1I4620_DIB[14], _6I4614_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_412_13 (_6I4614_$1I4488_$1I4620_DIB[13], _6I4614_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_412_12 (_6I4614_$1I4488_$1I4620_DIB[12], _6I4614_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_412_11 (_6I4614_$1I4488_$1I4620_DIB[11], _6I4614_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_412_10 (_6I4614_$1I4488_$1I4620_DIB[10], _6I4614_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_412_9 (_6I4614_$1I4488_$1I4620_DIB[9], _6I4614_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_412_8 (_6I4614_$1I4488_$1I4620_DIB[8], _6I4614_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_412_7 (_6I4614_$1I4488_$1I4620_DIB[7], _6I4614_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_412_6 (_6I4614_$1I4488_$1I4620_DIB[6], _6I4614_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_412_5 (_6I4614_$1I4488_$1I4620_DIB[5], _6I4614_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_412_4 (_6I4614_$1I4488_$1I4620_DIB[4], _6I4614_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_412_3 (_6I4614_$1I4488_$1I4620_DIB[3], _6I4614_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_412_2 (_6I4614_$1I4488_$1I4620_DIB[2], _6I4614_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_412_1 (_6I4614_$1I4488_$1I4620_DIB[1], _6I4614_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_412_0 (_6I4614_$1I4488_$1I4620_DIB[0], _6I4614_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _6I4614_$1I4488_$1I4620_DIPA;
 reg [1:16] _6I4614_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_413_0 (_6I4614_$1I4488_$1I4620_DIPA[0], _6I4614_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _6I4614_$1I4488_$1I4620_DIPB;
 reg [1:16] _6I4614_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_414_1 (_6I4614_$1I4488_$1I4620_DIPB[1], _6I4614_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _6I4614_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_414_0 (_6I4614_$1I4488_$1I4620_DIPB[0], _6I4614_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _6I4614_$1I4488_$1I4620_ENA;
 reg [1:16] _6I4614_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_415 (_6I4614_$1I4488_$1I4620_ENA, _6I4614_$1I4488_$1I4620_ENA__vlIN);

 wire  _6I4614_$1I4488_$1I4620_ENB;
 reg [1:16] _6I4614_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_416 (_6I4614_$1I4488_$1I4620_ENB, _6I4614_$1I4488_$1I4620_ENB__vlIN);

 wire  _6I4614_$1I4488_$1I4620_SSRA;
 reg [1:16] _6I4614_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_417 (_6I4614_$1I4488_$1I4620_SSRA, _6I4614_$1I4488_$1I4620_SSRA__vlIN);

 wire  _6I4614_$1I4488_$1I4620_SSRB;
 reg [1:16] _6I4614_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_418 (_6I4614_$1I4488_$1I4620_SSRB, _6I4614_$1I4488_$1I4620_SSRB__vlIN);

 wire  _6I4614_$1I4488_$1I4620_WEA;
 reg [1:16] _6I4614_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_419 (_6I4614_$1I4488_$1I4620_WEA, _6I4614_$1I4488_$1I4620_WEA__vlIN);

 wire  _6I4614_$1I4488_$1I4620_WEB;
 reg [1:16] _6I4614_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_420 (_6I4614_$1I4488_$1I4620_WEB, _6I4614_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _6I4614_$1I4488_$1I4620 ( _6I4614_$1I4488_$1I4620_DOA , _6I4614_$1I4488_$1I4620_DOB , _6I4614_$1I4488_$1I4620_DOPA , _6I4614_$1I4488_$1I4620_DOPB , _6I4614_$1I4488_$1I4620_ADDRA , _6I4614_$1I4488_$1I4620_ADDRB , _6I4614_$1I4488_$1I4620_CLKA , _6I4614_$1I4488_$1I4620_CLKB , _6I4614_$1I4488_$1I4620_DIA , _6I4614_$1I4488_$1I4620_DIB , _6I4614_$1I4488_$1I4620_DIPA , _6I4614_$1I4488_$1I4620_DIPB , _6I4614_$1I4488_$1I4620_ENA , _6I4614_$1I4488_$1I4620_ENB , _6I4614_$1I4488_$1I4620_SSRA , _6I4614_$1I4488_$1I4620_SSRB , _6I4614_$1I4488_$1I4620_WEA , _6I4614_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4598_$1I4488_$1I4621_DOA;

 wire [15:0] _6I4598_$1I4488_$1I4621_DOB;

 wire [0:0] _6I4598_$1I4488_$1I4621_DOPA;

 wire [1:0] _6I4598_$1I4488_$1I4621_DOPB;

 wire [10:0] _6I4598_$1I4488_$1I4621_ADDRA;
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_421_10 (_6I4598_$1I4488_$1I4621_ADDRA[10], _6I4598_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_421_9 (_6I4598_$1I4488_$1I4621_ADDRA[9], _6I4598_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_421_8 (_6I4598_$1I4488_$1I4621_ADDRA[8], _6I4598_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_421_7 (_6I4598_$1I4488_$1I4621_ADDRA[7], _6I4598_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_421_6 (_6I4598_$1I4488_$1I4621_ADDRA[6], _6I4598_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_421_5 (_6I4598_$1I4488_$1I4621_ADDRA[5], _6I4598_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_421_4 (_6I4598_$1I4488_$1I4621_ADDRA[4], _6I4598_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_421_3 (_6I4598_$1I4488_$1I4621_ADDRA[3], _6I4598_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_421_2 (_6I4598_$1I4488_$1I4621_ADDRA[2], _6I4598_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_421_1 (_6I4598_$1I4488_$1I4621_ADDRA[1], _6I4598_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_421_0 (_6I4598_$1I4488_$1I4621_ADDRA[0], _6I4598_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _6I4598_$1I4488_$1I4621_ADDRB;
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_422_9 (_6I4598_$1I4488_$1I4621_ADDRB[9], _6I4598_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_422_8 (_6I4598_$1I4488_$1I4621_ADDRB[8], _6I4598_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_422_7 (_6I4598_$1I4488_$1I4621_ADDRB[7], _6I4598_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_422_6 (_6I4598_$1I4488_$1I4621_ADDRB[6], _6I4598_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_422_5 (_6I4598_$1I4488_$1I4621_ADDRB[5], _6I4598_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_422_4 (_6I4598_$1I4488_$1I4621_ADDRB[4], _6I4598_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_422_3 (_6I4598_$1I4488_$1I4621_ADDRB[3], _6I4598_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_422_2 (_6I4598_$1I4488_$1I4621_ADDRB[2], _6I4598_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_422_1 (_6I4598_$1I4488_$1I4621_ADDRB[1], _6I4598_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_422_0 (_6I4598_$1I4488_$1I4621_ADDRB[0], _6I4598_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _6I4598_$1I4488_$1I4621_CLKA;
 reg [1:16] _6I4598_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_423 (_6I4598_$1I4488_$1I4621_CLKA, _6I4598_$1I4488_$1I4621_CLKA__vlIN);

 wire  _6I4598_$1I4488_$1I4621_CLKB;
 reg [1:16] _6I4598_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_424 (_6I4598_$1I4488_$1I4621_CLKB, _6I4598_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _6I4598_$1I4488_$1I4621_DIA;
 reg [1:16] _6I4598_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_425_7 (_6I4598_$1I4488_$1I4621_DIA[7], _6I4598_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_425_6 (_6I4598_$1I4488_$1I4621_DIA[6], _6I4598_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_425_5 (_6I4598_$1I4488_$1I4621_DIA[5], _6I4598_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_425_4 (_6I4598_$1I4488_$1I4621_DIA[4], _6I4598_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_425_3 (_6I4598_$1I4488_$1I4621_DIA[3], _6I4598_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_425_2 (_6I4598_$1I4488_$1I4621_DIA[2], _6I4598_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_425_1 (_6I4598_$1I4488_$1I4621_DIA[1], _6I4598_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_425_0 (_6I4598_$1I4488_$1I4621_DIA[0], _6I4598_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _6I4598_$1I4488_$1I4621_DIB;
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_426_15 (_6I4598_$1I4488_$1I4621_DIB[15], _6I4598_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_426_14 (_6I4598_$1I4488_$1I4621_DIB[14], _6I4598_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_426_13 (_6I4598_$1I4488_$1I4621_DIB[13], _6I4598_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_426_12 (_6I4598_$1I4488_$1I4621_DIB[12], _6I4598_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_426_11 (_6I4598_$1I4488_$1I4621_DIB[11], _6I4598_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_426_10 (_6I4598_$1I4488_$1I4621_DIB[10], _6I4598_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_426_9 (_6I4598_$1I4488_$1I4621_DIB[9], _6I4598_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_426_8 (_6I4598_$1I4488_$1I4621_DIB[8], _6I4598_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_426_7 (_6I4598_$1I4488_$1I4621_DIB[7], _6I4598_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_426_6 (_6I4598_$1I4488_$1I4621_DIB[6], _6I4598_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_426_5 (_6I4598_$1I4488_$1I4621_DIB[5], _6I4598_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_426_4 (_6I4598_$1I4488_$1I4621_DIB[4], _6I4598_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_426_3 (_6I4598_$1I4488_$1I4621_DIB[3], _6I4598_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_426_2 (_6I4598_$1I4488_$1I4621_DIB[2], _6I4598_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_426_1 (_6I4598_$1I4488_$1I4621_DIB[1], _6I4598_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_426_0 (_6I4598_$1I4488_$1I4621_DIB[0], _6I4598_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _6I4598_$1I4488_$1I4621_DIPA;
 reg [1:16] _6I4598_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_427_0 (_6I4598_$1I4488_$1I4621_DIPA[0], _6I4598_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _6I4598_$1I4488_$1I4621_DIPB;
 reg [1:16] _6I4598_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_428_1 (_6I4598_$1I4488_$1I4621_DIPB[1], _6I4598_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_428_0 (_6I4598_$1I4488_$1I4621_DIPB[0], _6I4598_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _6I4598_$1I4488_$1I4621_ENA;
 reg [1:16] _6I4598_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_429 (_6I4598_$1I4488_$1I4621_ENA, _6I4598_$1I4488_$1I4621_ENA__vlIN);

 wire  _6I4598_$1I4488_$1I4621_ENB;
 reg [1:16] _6I4598_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_430 (_6I4598_$1I4488_$1I4621_ENB, _6I4598_$1I4488_$1I4621_ENB__vlIN);

 wire  _6I4598_$1I4488_$1I4621_SSRA;
 reg [1:16] _6I4598_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_431 (_6I4598_$1I4488_$1I4621_SSRA, _6I4598_$1I4488_$1I4621_SSRA__vlIN);

 wire  _6I4598_$1I4488_$1I4621_SSRB;
 reg [1:16] _6I4598_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_432 (_6I4598_$1I4488_$1I4621_SSRB, _6I4598_$1I4488_$1I4621_SSRB__vlIN);

 wire  _6I4598_$1I4488_$1I4621_WEA;
 reg [1:16] _6I4598_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_433 (_6I4598_$1I4488_$1I4621_WEA, _6I4598_$1I4488_$1I4621_WEA__vlIN);

 wire  _6I4598_$1I4488_$1I4621_WEB;
 reg [1:16] _6I4598_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_434 (_6I4598_$1I4488_$1I4621_WEB, _6I4598_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _6I4598_$1I4488_$1I4621 ( _6I4598_$1I4488_$1I4621_DOA , _6I4598_$1I4488_$1I4621_DOB , _6I4598_$1I4488_$1I4621_DOPA , _6I4598_$1I4488_$1I4621_DOPB , _6I4598_$1I4488_$1I4621_ADDRA , _6I4598_$1I4488_$1I4621_ADDRB , _6I4598_$1I4488_$1I4621_CLKA , _6I4598_$1I4488_$1I4621_CLKB , _6I4598_$1I4488_$1I4621_DIA , _6I4598_$1I4488_$1I4621_DIB , _6I4598_$1I4488_$1I4621_DIPA , _6I4598_$1I4488_$1I4621_DIPB , _6I4598_$1I4488_$1I4621_ENA , _6I4598_$1I4488_$1I4621_ENB , _6I4598_$1I4488_$1I4621_SSRA , _6I4598_$1I4488_$1I4621_SSRB , _6I4598_$1I4488_$1I4621_WEA , _6I4598_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4598_$1I4488_$1I4620_DOA;

 wire [15:0] _6I4598_$1I4488_$1I4620_DOB;

 wire [0:0] _6I4598_$1I4488_$1I4620_DOPA;

 wire [1:0] _6I4598_$1I4488_$1I4620_DOPB;

 wire [10:0] _6I4598_$1I4488_$1I4620_ADDRA;
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_435_10 (_6I4598_$1I4488_$1I4620_ADDRA[10], _6I4598_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_435_9 (_6I4598_$1I4488_$1I4620_ADDRA[9], _6I4598_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_435_8 (_6I4598_$1I4488_$1I4620_ADDRA[8], _6I4598_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_435_7 (_6I4598_$1I4488_$1I4620_ADDRA[7], _6I4598_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_435_6 (_6I4598_$1I4488_$1I4620_ADDRA[6], _6I4598_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_435_5 (_6I4598_$1I4488_$1I4620_ADDRA[5], _6I4598_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_435_4 (_6I4598_$1I4488_$1I4620_ADDRA[4], _6I4598_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_435_3 (_6I4598_$1I4488_$1I4620_ADDRA[3], _6I4598_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_435_2 (_6I4598_$1I4488_$1I4620_ADDRA[2], _6I4598_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_435_1 (_6I4598_$1I4488_$1I4620_ADDRA[1], _6I4598_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_435_0 (_6I4598_$1I4488_$1I4620_ADDRA[0], _6I4598_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _6I4598_$1I4488_$1I4620_ADDRB;
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_436_9 (_6I4598_$1I4488_$1I4620_ADDRB[9], _6I4598_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_436_8 (_6I4598_$1I4488_$1I4620_ADDRB[8], _6I4598_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_436_7 (_6I4598_$1I4488_$1I4620_ADDRB[7], _6I4598_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_436_6 (_6I4598_$1I4488_$1I4620_ADDRB[6], _6I4598_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_436_5 (_6I4598_$1I4488_$1I4620_ADDRB[5], _6I4598_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_436_4 (_6I4598_$1I4488_$1I4620_ADDRB[4], _6I4598_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_436_3 (_6I4598_$1I4488_$1I4620_ADDRB[3], _6I4598_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_436_2 (_6I4598_$1I4488_$1I4620_ADDRB[2], _6I4598_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_436_1 (_6I4598_$1I4488_$1I4620_ADDRB[1], _6I4598_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_436_0 (_6I4598_$1I4488_$1I4620_ADDRB[0], _6I4598_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _6I4598_$1I4488_$1I4620_CLKA;
 reg [1:16] _6I4598_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_437 (_6I4598_$1I4488_$1I4620_CLKA, _6I4598_$1I4488_$1I4620_CLKA__vlIN);

 wire  _6I4598_$1I4488_$1I4620_CLKB;
 reg [1:16] _6I4598_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_438 (_6I4598_$1I4488_$1I4620_CLKB, _6I4598_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _6I4598_$1I4488_$1I4620_DIA;
 reg [1:16] _6I4598_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_439_7 (_6I4598_$1I4488_$1I4620_DIA[7], _6I4598_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_439_6 (_6I4598_$1I4488_$1I4620_DIA[6], _6I4598_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_439_5 (_6I4598_$1I4488_$1I4620_DIA[5], _6I4598_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_439_4 (_6I4598_$1I4488_$1I4620_DIA[4], _6I4598_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_439_3 (_6I4598_$1I4488_$1I4620_DIA[3], _6I4598_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_439_2 (_6I4598_$1I4488_$1I4620_DIA[2], _6I4598_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_439_1 (_6I4598_$1I4488_$1I4620_DIA[1], _6I4598_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_439_0 (_6I4598_$1I4488_$1I4620_DIA[0], _6I4598_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _6I4598_$1I4488_$1I4620_DIB;
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_440_15 (_6I4598_$1I4488_$1I4620_DIB[15], _6I4598_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_440_14 (_6I4598_$1I4488_$1I4620_DIB[14], _6I4598_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_440_13 (_6I4598_$1I4488_$1I4620_DIB[13], _6I4598_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_440_12 (_6I4598_$1I4488_$1I4620_DIB[12], _6I4598_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_440_11 (_6I4598_$1I4488_$1I4620_DIB[11], _6I4598_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_440_10 (_6I4598_$1I4488_$1I4620_DIB[10], _6I4598_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_440_9 (_6I4598_$1I4488_$1I4620_DIB[9], _6I4598_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_440_8 (_6I4598_$1I4488_$1I4620_DIB[8], _6I4598_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_440_7 (_6I4598_$1I4488_$1I4620_DIB[7], _6I4598_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_440_6 (_6I4598_$1I4488_$1I4620_DIB[6], _6I4598_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_440_5 (_6I4598_$1I4488_$1I4620_DIB[5], _6I4598_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_440_4 (_6I4598_$1I4488_$1I4620_DIB[4], _6I4598_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_440_3 (_6I4598_$1I4488_$1I4620_DIB[3], _6I4598_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_440_2 (_6I4598_$1I4488_$1I4620_DIB[2], _6I4598_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_440_1 (_6I4598_$1I4488_$1I4620_DIB[1], _6I4598_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_440_0 (_6I4598_$1I4488_$1I4620_DIB[0], _6I4598_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _6I4598_$1I4488_$1I4620_DIPA;
 reg [1:16] _6I4598_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_441_0 (_6I4598_$1I4488_$1I4620_DIPA[0], _6I4598_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _6I4598_$1I4488_$1I4620_DIPB;
 reg [1:16] _6I4598_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_442_1 (_6I4598_$1I4488_$1I4620_DIPB[1], _6I4598_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _6I4598_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_442_0 (_6I4598_$1I4488_$1I4620_DIPB[0], _6I4598_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _6I4598_$1I4488_$1I4620_ENA;
 reg [1:16] _6I4598_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_443 (_6I4598_$1I4488_$1I4620_ENA, _6I4598_$1I4488_$1I4620_ENA__vlIN);

 wire  _6I4598_$1I4488_$1I4620_ENB;
 reg [1:16] _6I4598_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_444 (_6I4598_$1I4488_$1I4620_ENB, _6I4598_$1I4488_$1I4620_ENB__vlIN);

 wire  _6I4598_$1I4488_$1I4620_SSRA;
 reg [1:16] _6I4598_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_445 (_6I4598_$1I4488_$1I4620_SSRA, _6I4598_$1I4488_$1I4620_SSRA__vlIN);

 wire  _6I4598_$1I4488_$1I4620_SSRB;
 reg [1:16] _6I4598_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_446 (_6I4598_$1I4488_$1I4620_SSRB, _6I4598_$1I4488_$1I4620_SSRB__vlIN);

 wire  _6I4598_$1I4488_$1I4620_WEA;
 reg [1:16] _6I4598_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_447 (_6I4598_$1I4488_$1I4620_WEA, _6I4598_$1I4488_$1I4620_WEA__vlIN);

 wire  _6I4598_$1I4488_$1I4620_WEB;
 reg [1:16] _6I4598_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_448 (_6I4598_$1I4488_$1I4620_WEB, _6I4598_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _6I4598_$1I4488_$1I4620 ( _6I4598_$1I4488_$1I4620_DOA , _6I4598_$1I4488_$1I4620_DOB , _6I4598_$1I4488_$1I4620_DOPA , _6I4598_$1I4488_$1I4620_DOPB , _6I4598_$1I4488_$1I4620_ADDRA , _6I4598_$1I4488_$1I4620_ADDRB , _6I4598_$1I4488_$1I4620_CLKA , _6I4598_$1I4488_$1I4620_CLKB , _6I4598_$1I4488_$1I4620_DIA , _6I4598_$1I4488_$1I4620_DIB , _6I4598_$1I4488_$1I4620_DIPA , _6I4598_$1I4488_$1I4620_DIPB , _6I4598_$1I4488_$1I4620_ENA , _6I4598_$1I4488_$1I4620_ENB , _6I4598_$1I4488_$1I4620_SSRA , _6I4598_$1I4488_$1I4620_SSRB , _6I4598_$1I4488_$1I4620_WEA , _6I4598_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4575_$1I4488_$1I4621_DOA;

 wire [15:0] _6I4575_$1I4488_$1I4621_DOB;

 wire [0:0] _6I4575_$1I4488_$1I4621_DOPA;

 wire [1:0] _6I4575_$1I4488_$1I4621_DOPB;

 wire [10:0] _6I4575_$1I4488_$1I4621_ADDRA;
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_449_10 (_6I4575_$1I4488_$1I4621_ADDRA[10], _6I4575_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_449_9 (_6I4575_$1I4488_$1I4621_ADDRA[9], _6I4575_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_449_8 (_6I4575_$1I4488_$1I4621_ADDRA[8], _6I4575_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_449_7 (_6I4575_$1I4488_$1I4621_ADDRA[7], _6I4575_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_449_6 (_6I4575_$1I4488_$1I4621_ADDRA[6], _6I4575_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_449_5 (_6I4575_$1I4488_$1I4621_ADDRA[5], _6I4575_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_449_4 (_6I4575_$1I4488_$1I4621_ADDRA[4], _6I4575_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_449_3 (_6I4575_$1I4488_$1I4621_ADDRA[3], _6I4575_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_449_2 (_6I4575_$1I4488_$1I4621_ADDRA[2], _6I4575_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_449_1 (_6I4575_$1I4488_$1I4621_ADDRA[1], _6I4575_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_449_0 (_6I4575_$1I4488_$1I4621_ADDRA[0], _6I4575_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _6I4575_$1I4488_$1I4621_ADDRB;
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_450_9 (_6I4575_$1I4488_$1I4621_ADDRB[9], _6I4575_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_450_8 (_6I4575_$1I4488_$1I4621_ADDRB[8], _6I4575_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_450_7 (_6I4575_$1I4488_$1I4621_ADDRB[7], _6I4575_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_450_6 (_6I4575_$1I4488_$1I4621_ADDRB[6], _6I4575_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_450_5 (_6I4575_$1I4488_$1I4621_ADDRB[5], _6I4575_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_450_4 (_6I4575_$1I4488_$1I4621_ADDRB[4], _6I4575_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_450_3 (_6I4575_$1I4488_$1I4621_ADDRB[3], _6I4575_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_450_2 (_6I4575_$1I4488_$1I4621_ADDRB[2], _6I4575_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_450_1 (_6I4575_$1I4488_$1I4621_ADDRB[1], _6I4575_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_450_0 (_6I4575_$1I4488_$1I4621_ADDRB[0], _6I4575_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _6I4575_$1I4488_$1I4621_CLKA;
 reg [1:16] _6I4575_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_451 (_6I4575_$1I4488_$1I4621_CLKA, _6I4575_$1I4488_$1I4621_CLKA__vlIN);

 wire  _6I4575_$1I4488_$1I4621_CLKB;
 reg [1:16] _6I4575_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_452 (_6I4575_$1I4488_$1I4621_CLKB, _6I4575_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _6I4575_$1I4488_$1I4621_DIA;
 reg [1:16] _6I4575_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_453_7 (_6I4575_$1I4488_$1I4621_DIA[7], _6I4575_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_453_6 (_6I4575_$1I4488_$1I4621_DIA[6], _6I4575_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_453_5 (_6I4575_$1I4488_$1I4621_DIA[5], _6I4575_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_453_4 (_6I4575_$1I4488_$1I4621_DIA[4], _6I4575_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_453_3 (_6I4575_$1I4488_$1I4621_DIA[3], _6I4575_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_453_2 (_6I4575_$1I4488_$1I4621_DIA[2], _6I4575_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_453_1 (_6I4575_$1I4488_$1I4621_DIA[1], _6I4575_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_453_0 (_6I4575_$1I4488_$1I4621_DIA[0], _6I4575_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _6I4575_$1I4488_$1I4621_DIB;
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_454_15 (_6I4575_$1I4488_$1I4621_DIB[15], _6I4575_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_454_14 (_6I4575_$1I4488_$1I4621_DIB[14], _6I4575_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_454_13 (_6I4575_$1I4488_$1I4621_DIB[13], _6I4575_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_454_12 (_6I4575_$1I4488_$1I4621_DIB[12], _6I4575_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_454_11 (_6I4575_$1I4488_$1I4621_DIB[11], _6I4575_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_454_10 (_6I4575_$1I4488_$1I4621_DIB[10], _6I4575_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_454_9 (_6I4575_$1I4488_$1I4621_DIB[9], _6I4575_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_454_8 (_6I4575_$1I4488_$1I4621_DIB[8], _6I4575_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_454_7 (_6I4575_$1I4488_$1I4621_DIB[7], _6I4575_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_454_6 (_6I4575_$1I4488_$1I4621_DIB[6], _6I4575_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_454_5 (_6I4575_$1I4488_$1I4621_DIB[5], _6I4575_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_454_4 (_6I4575_$1I4488_$1I4621_DIB[4], _6I4575_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_454_3 (_6I4575_$1I4488_$1I4621_DIB[3], _6I4575_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_454_2 (_6I4575_$1I4488_$1I4621_DIB[2], _6I4575_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_454_1 (_6I4575_$1I4488_$1I4621_DIB[1], _6I4575_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_454_0 (_6I4575_$1I4488_$1I4621_DIB[0], _6I4575_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _6I4575_$1I4488_$1I4621_DIPA;
 reg [1:16] _6I4575_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_455_0 (_6I4575_$1I4488_$1I4621_DIPA[0], _6I4575_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _6I4575_$1I4488_$1I4621_DIPB;
 reg [1:16] _6I4575_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_456_1 (_6I4575_$1I4488_$1I4621_DIPB[1], _6I4575_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_456_0 (_6I4575_$1I4488_$1I4621_DIPB[0], _6I4575_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _6I4575_$1I4488_$1I4621_ENA;
 reg [1:16] _6I4575_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_457 (_6I4575_$1I4488_$1I4621_ENA, _6I4575_$1I4488_$1I4621_ENA__vlIN);

 wire  _6I4575_$1I4488_$1I4621_ENB;
 reg [1:16] _6I4575_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_458 (_6I4575_$1I4488_$1I4621_ENB, _6I4575_$1I4488_$1I4621_ENB__vlIN);

 wire  _6I4575_$1I4488_$1I4621_SSRA;
 reg [1:16] _6I4575_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_459 (_6I4575_$1I4488_$1I4621_SSRA, _6I4575_$1I4488_$1I4621_SSRA__vlIN);

 wire  _6I4575_$1I4488_$1I4621_SSRB;
 reg [1:16] _6I4575_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_460 (_6I4575_$1I4488_$1I4621_SSRB, _6I4575_$1I4488_$1I4621_SSRB__vlIN);

 wire  _6I4575_$1I4488_$1I4621_WEA;
 reg [1:16] _6I4575_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_461 (_6I4575_$1I4488_$1I4621_WEA, _6I4575_$1I4488_$1I4621_WEA__vlIN);

 wire  _6I4575_$1I4488_$1I4621_WEB;
 reg [1:16] _6I4575_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_462 (_6I4575_$1I4488_$1I4621_WEB, _6I4575_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _6I4575_$1I4488_$1I4621 ( _6I4575_$1I4488_$1I4621_DOA , _6I4575_$1I4488_$1I4621_DOB , _6I4575_$1I4488_$1I4621_DOPA , _6I4575_$1I4488_$1I4621_DOPB , _6I4575_$1I4488_$1I4621_ADDRA , _6I4575_$1I4488_$1I4621_ADDRB , _6I4575_$1I4488_$1I4621_CLKA , _6I4575_$1I4488_$1I4621_CLKB , _6I4575_$1I4488_$1I4621_DIA , _6I4575_$1I4488_$1I4621_DIB , _6I4575_$1I4488_$1I4621_DIPA , _6I4575_$1I4488_$1I4621_DIPB , _6I4575_$1I4488_$1I4621_ENA , _6I4575_$1I4488_$1I4621_ENB , _6I4575_$1I4488_$1I4621_SSRA , _6I4575_$1I4488_$1I4621_SSRB , _6I4575_$1I4488_$1I4621_WEA , _6I4575_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4575_$1I4488_$1I4620_DOA;

 wire [15:0] _6I4575_$1I4488_$1I4620_DOB;

 wire [0:0] _6I4575_$1I4488_$1I4620_DOPA;

 wire [1:0] _6I4575_$1I4488_$1I4620_DOPB;

 wire [10:0] _6I4575_$1I4488_$1I4620_ADDRA;
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_463_10 (_6I4575_$1I4488_$1I4620_ADDRA[10], _6I4575_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_463_9 (_6I4575_$1I4488_$1I4620_ADDRA[9], _6I4575_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_463_8 (_6I4575_$1I4488_$1I4620_ADDRA[8], _6I4575_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_463_7 (_6I4575_$1I4488_$1I4620_ADDRA[7], _6I4575_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_463_6 (_6I4575_$1I4488_$1I4620_ADDRA[6], _6I4575_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_463_5 (_6I4575_$1I4488_$1I4620_ADDRA[5], _6I4575_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_463_4 (_6I4575_$1I4488_$1I4620_ADDRA[4], _6I4575_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_463_3 (_6I4575_$1I4488_$1I4620_ADDRA[3], _6I4575_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_463_2 (_6I4575_$1I4488_$1I4620_ADDRA[2], _6I4575_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_463_1 (_6I4575_$1I4488_$1I4620_ADDRA[1], _6I4575_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_463_0 (_6I4575_$1I4488_$1I4620_ADDRA[0], _6I4575_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _6I4575_$1I4488_$1I4620_ADDRB;
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_464_9 (_6I4575_$1I4488_$1I4620_ADDRB[9], _6I4575_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_464_8 (_6I4575_$1I4488_$1I4620_ADDRB[8], _6I4575_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_464_7 (_6I4575_$1I4488_$1I4620_ADDRB[7], _6I4575_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_464_6 (_6I4575_$1I4488_$1I4620_ADDRB[6], _6I4575_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_464_5 (_6I4575_$1I4488_$1I4620_ADDRB[5], _6I4575_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_464_4 (_6I4575_$1I4488_$1I4620_ADDRB[4], _6I4575_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_464_3 (_6I4575_$1I4488_$1I4620_ADDRB[3], _6I4575_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_464_2 (_6I4575_$1I4488_$1I4620_ADDRB[2], _6I4575_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_464_1 (_6I4575_$1I4488_$1I4620_ADDRB[1], _6I4575_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_464_0 (_6I4575_$1I4488_$1I4620_ADDRB[0], _6I4575_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _6I4575_$1I4488_$1I4620_CLKA;
 reg [1:16] _6I4575_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_465 (_6I4575_$1I4488_$1I4620_CLKA, _6I4575_$1I4488_$1I4620_CLKA__vlIN);

 wire  _6I4575_$1I4488_$1I4620_CLKB;
 reg [1:16] _6I4575_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_466 (_6I4575_$1I4488_$1I4620_CLKB, _6I4575_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _6I4575_$1I4488_$1I4620_DIA;
 reg [1:16] _6I4575_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_467_7 (_6I4575_$1I4488_$1I4620_DIA[7], _6I4575_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_467_6 (_6I4575_$1I4488_$1I4620_DIA[6], _6I4575_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_467_5 (_6I4575_$1I4488_$1I4620_DIA[5], _6I4575_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_467_4 (_6I4575_$1I4488_$1I4620_DIA[4], _6I4575_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_467_3 (_6I4575_$1I4488_$1I4620_DIA[3], _6I4575_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_467_2 (_6I4575_$1I4488_$1I4620_DIA[2], _6I4575_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_467_1 (_6I4575_$1I4488_$1I4620_DIA[1], _6I4575_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_467_0 (_6I4575_$1I4488_$1I4620_DIA[0], _6I4575_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _6I4575_$1I4488_$1I4620_DIB;
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_468_15 (_6I4575_$1I4488_$1I4620_DIB[15], _6I4575_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_468_14 (_6I4575_$1I4488_$1I4620_DIB[14], _6I4575_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_468_13 (_6I4575_$1I4488_$1I4620_DIB[13], _6I4575_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_468_12 (_6I4575_$1I4488_$1I4620_DIB[12], _6I4575_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_468_11 (_6I4575_$1I4488_$1I4620_DIB[11], _6I4575_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_468_10 (_6I4575_$1I4488_$1I4620_DIB[10], _6I4575_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_468_9 (_6I4575_$1I4488_$1I4620_DIB[9], _6I4575_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_468_8 (_6I4575_$1I4488_$1I4620_DIB[8], _6I4575_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_468_7 (_6I4575_$1I4488_$1I4620_DIB[7], _6I4575_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_468_6 (_6I4575_$1I4488_$1I4620_DIB[6], _6I4575_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_468_5 (_6I4575_$1I4488_$1I4620_DIB[5], _6I4575_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_468_4 (_6I4575_$1I4488_$1I4620_DIB[4], _6I4575_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_468_3 (_6I4575_$1I4488_$1I4620_DIB[3], _6I4575_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_468_2 (_6I4575_$1I4488_$1I4620_DIB[2], _6I4575_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_468_1 (_6I4575_$1I4488_$1I4620_DIB[1], _6I4575_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_468_0 (_6I4575_$1I4488_$1I4620_DIB[0], _6I4575_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _6I4575_$1I4488_$1I4620_DIPA;
 reg [1:16] _6I4575_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_469_0 (_6I4575_$1I4488_$1I4620_DIPA[0], _6I4575_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _6I4575_$1I4488_$1I4620_DIPB;
 reg [1:16] _6I4575_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_470_1 (_6I4575_$1I4488_$1I4620_DIPB[1], _6I4575_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _6I4575_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_470_0 (_6I4575_$1I4488_$1I4620_DIPB[0], _6I4575_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _6I4575_$1I4488_$1I4620_ENA;
 reg [1:16] _6I4575_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_471 (_6I4575_$1I4488_$1I4620_ENA, _6I4575_$1I4488_$1I4620_ENA__vlIN);

 wire  _6I4575_$1I4488_$1I4620_ENB;
 reg [1:16] _6I4575_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_472 (_6I4575_$1I4488_$1I4620_ENB, _6I4575_$1I4488_$1I4620_ENB__vlIN);

 wire  _6I4575_$1I4488_$1I4620_SSRA;
 reg [1:16] _6I4575_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_473 (_6I4575_$1I4488_$1I4620_SSRA, _6I4575_$1I4488_$1I4620_SSRA__vlIN);

 wire  _6I4575_$1I4488_$1I4620_SSRB;
 reg [1:16] _6I4575_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_474 (_6I4575_$1I4488_$1I4620_SSRB, _6I4575_$1I4488_$1I4620_SSRB__vlIN);

 wire  _6I4575_$1I4488_$1I4620_WEA;
 reg [1:16] _6I4575_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_475 (_6I4575_$1I4488_$1I4620_WEA, _6I4575_$1I4488_$1I4620_WEA__vlIN);

 wire  _6I4575_$1I4488_$1I4620_WEB;
 reg [1:16] _6I4575_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_476 (_6I4575_$1I4488_$1I4620_WEB, _6I4575_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _6I4575_$1I4488_$1I4620 ( _6I4575_$1I4488_$1I4620_DOA , _6I4575_$1I4488_$1I4620_DOB , _6I4575_$1I4488_$1I4620_DOPA , _6I4575_$1I4488_$1I4620_DOPB , _6I4575_$1I4488_$1I4620_ADDRA , _6I4575_$1I4488_$1I4620_ADDRB , _6I4575_$1I4488_$1I4620_CLKA , _6I4575_$1I4488_$1I4620_CLKB , _6I4575_$1I4488_$1I4620_DIA , _6I4575_$1I4488_$1I4620_DIB , _6I4575_$1I4488_$1I4620_DIPA , _6I4575_$1I4488_$1I4620_DIPB , _6I4575_$1I4488_$1I4620_ENA , _6I4575_$1I4488_$1I4620_ENB , _6I4575_$1I4488_$1I4620_SSRA , _6I4575_$1I4488_$1I4620_SSRB , _6I4575_$1I4488_$1I4620_WEA , _6I4575_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4529_$1I4488_$1I4621_DOA;

 wire [15:0] _6I4529_$1I4488_$1I4621_DOB;

 wire [0:0] _6I4529_$1I4488_$1I4621_DOPA;

 wire [1:0] _6I4529_$1I4488_$1I4621_DOPB;

 wire [10:0] _6I4529_$1I4488_$1I4621_ADDRA;
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_477_10 (_6I4529_$1I4488_$1I4621_ADDRA[10], _6I4529_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_477_9 (_6I4529_$1I4488_$1I4621_ADDRA[9], _6I4529_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_477_8 (_6I4529_$1I4488_$1I4621_ADDRA[8], _6I4529_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_477_7 (_6I4529_$1I4488_$1I4621_ADDRA[7], _6I4529_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_477_6 (_6I4529_$1I4488_$1I4621_ADDRA[6], _6I4529_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_477_5 (_6I4529_$1I4488_$1I4621_ADDRA[5], _6I4529_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_477_4 (_6I4529_$1I4488_$1I4621_ADDRA[4], _6I4529_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_477_3 (_6I4529_$1I4488_$1I4621_ADDRA[3], _6I4529_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_477_2 (_6I4529_$1I4488_$1I4621_ADDRA[2], _6I4529_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_477_1 (_6I4529_$1I4488_$1I4621_ADDRA[1], _6I4529_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_477_0 (_6I4529_$1I4488_$1I4621_ADDRA[0], _6I4529_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _6I4529_$1I4488_$1I4621_ADDRB;
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_478_9 (_6I4529_$1I4488_$1I4621_ADDRB[9], _6I4529_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_478_8 (_6I4529_$1I4488_$1I4621_ADDRB[8], _6I4529_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_478_7 (_6I4529_$1I4488_$1I4621_ADDRB[7], _6I4529_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_478_6 (_6I4529_$1I4488_$1I4621_ADDRB[6], _6I4529_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_478_5 (_6I4529_$1I4488_$1I4621_ADDRB[5], _6I4529_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_478_4 (_6I4529_$1I4488_$1I4621_ADDRB[4], _6I4529_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_478_3 (_6I4529_$1I4488_$1I4621_ADDRB[3], _6I4529_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_478_2 (_6I4529_$1I4488_$1I4621_ADDRB[2], _6I4529_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_478_1 (_6I4529_$1I4488_$1I4621_ADDRB[1], _6I4529_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_478_0 (_6I4529_$1I4488_$1I4621_ADDRB[0], _6I4529_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _6I4529_$1I4488_$1I4621_CLKA;
 reg [1:16] _6I4529_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_479 (_6I4529_$1I4488_$1I4621_CLKA, _6I4529_$1I4488_$1I4621_CLKA__vlIN);

 wire  _6I4529_$1I4488_$1I4621_CLKB;
 reg [1:16] _6I4529_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_480 (_6I4529_$1I4488_$1I4621_CLKB, _6I4529_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _6I4529_$1I4488_$1I4621_DIA;
 reg [1:16] _6I4529_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_481_7 (_6I4529_$1I4488_$1I4621_DIA[7], _6I4529_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_481_6 (_6I4529_$1I4488_$1I4621_DIA[6], _6I4529_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_481_5 (_6I4529_$1I4488_$1I4621_DIA[5], _6I4529_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_481_4 (_6I4529_$1I4488_$1I4621_DIA[4], _6I4529_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_481_3 (_6I4529_$1I4488_$1I4621_DIA[3], _6I4529_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_481_2 (_6I4529_$1I4488_$1I4621_DIA[2], _6I4529_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_481_1 (_6I4529_$1I4488_$1I4621_DIA[1], _6I4529_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_481_0 (_6I4529_$1I4488_$1I4621_DIA[0], _6I4529_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _6I4529_$1I4488_$1I4621_DIB;
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_482_15 (_6I4529_$1I4488_$1I4621_DIB[15], _6I4529_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_482_14 (_6I4529_$1I4488_$1I4621_DIB[14], _6I4529_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_482_13 (_6I4529_$1I4488_$1I4621_DIB[13], _6I4529_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_482_12 (_6I4529_$1I4488_$1I4621_DIB[12], _6I4529_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_482_11 (_6I4529_$1I4488_$1I4621_DIB[11], _6I4529_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_482_10 (_6I4529_$1I4488_$1I4621_DIB[10], _6I4529_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_482_9 (_6I4529_$1I4488_$1I4621_DIB[9], _6I4529_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_482_8 (_6I4529_$1I4488_$1I4621_DIB[8], _6I4529_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_482_7 (_6I4529_$1I4488_$1I4621_DIB[7], _6I4529_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_482_6 (_6I4529_$1I4488_$1I4621_DIB[6], _6I4529_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_482_5 (_6I4529_$1I4488_$1I4621_DIB[5], _6I4529_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_482_4 (_6I4529_$1I4488_$1I4621_DIB[4], _6I4529_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_482_3 (_6I4529_$1I4488_$1I4621_DIB[3], _6I4529_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_482_2 (_6I4529_$1I4488_$1I4621_DIB[2], _6I4529_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_482_1 (_6I4529_$1I4488_$1I4621_DIB[1], _6I4529_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_482_0 (_6I4529_$1I4488_$1I4621_DIB[0], _6I4529_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _6I4529_$1I4488_$1I4621_DIPA;
 reg [1:16] _6I4529_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_483_0 (_6I4529_$1I4488_$1I4621_DIPA[0], _6I4529_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _6I4529_$1I4488_$1I4621_DIPB;
 reg [1:16] _6I4529_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_484_1 (_6I4529_$1I4488_$1I4621_DIPB[1], _6I4529_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_484_0 (_6I4529_$1I4488_$1I4621_DIPB[0], _6I4529_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _6I4529_$1I4488_$1I4621_ENA;
 reg [1:16] _6I4529_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_485 (_6I4529_$1I4488_$1I4621_ENA, _6I4529_$1I4488_$1I4621_ENA__vlIN);

 wire  _6I4529_$1I4488_$1I4621_ENB;
 reg [1:16] _6I4529_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_486 (_6I4529_$1I4488_$1I4621_ENB, _6I4529_$1I4488_$1I4621_ENB__vlIN);

 wire  _6I4529_$1I4488_$1I4621_SSRA;
 reg [1:16] _6I4529_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_487 (_6I4529_$1I4488_$1I4621_SSRA, _6I4529_$1I4488_$1I4621_SSRA__vlIN);

 wire  _6I4529_$1I4488_$1I4621_SSRB;
 reg [1:16] _6I4529_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_488 (_6I4529_$1I4488_$1I4621_SSRB, _6I4529_$1I4488_$1I4621_SSRB__vlIN);

 wire  _6I4529_$1I4488_$1I4621_WEA;
 reg [1:16] _6I4529_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_489 (_6I4529_$1I4488_$1I4621_WEA, _6I4529_$1I4488_$1I4621_WEA__vlIN);

 wire  _6I4529_$1I4488_$1I4621_WEB;
 reg [1:16] _6I4529_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_490 (_6I4529_$1I4488_$1I4621_WEB, _6I4529_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _6I4529_$1I4488_$1I4621 ( _6I4529_$1I4488_$1I4621_DOA , _6I4529_$1I4488_$1I4621_DOB , _6I4529_$1I4488_$1I4621_DOPA , _6I4529_$1I4488_$1I4621_DOPB , _6I4529_$1I4488_$1I4621_ADDRA , _6I4529_$1I4488_$1I4621_ADDRB , _6I4529_$1I4488_$1I4621_CLKA , _6I4529_$1I4488_$1I4621_CLKB , _6I4529_$1I4488_$1I4621_DIA , _6I4529_$1I4488_$1I4621_DIB , _6I4529_$1I4488_$1I4621_DIPA , _6I4529_$1I4488_$1I4621_DIPB , _6I4529_$1I4488_$1I4621_ENA , _6I4529_$1I4488_$1I4621_ENB , _6I4529_$1I4488_$1I4621_SSRA , _6I4529_$1I4488_$1I4621_SSRB , _6I4529_$1I4488_$1I4621_WEA , _6I4529_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4529_$1I4488_$1I4620_DOA;

 wire [15:0] _6I4529_$1I4488_$1I4620_DOB;

 wire [0:0] _6I4529_$1I4488_$1I4620_DOPA;

 wire [1:0] _6I4529_$1I4488_$1I4620_DOPB;

 wire [10:0] _6I4529_$1I4488_$1I4620_ADDRA;
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_491_10 (_6I4529_$1I4488_$1I4620_ADDRA[10], _6I4529_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_491_9 (_6I4529_$1I4488_$1I4620_ADDRA[9], _6I4529_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_491_8 (_6I4529_$1I4488_$1I4620_ADDRA[8], _6I4529_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_491_7 (_6I4529_$1I4488_$1I4620_ADDRA[7], _6I4529_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_491_6 (_6I4529_$1I4488_$1I4620_ADDRA[6], _6I4529_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_491_5 (_6I4529_$1I4488_$1I4620_ADDRA[5], _6I4529_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_491_4 (_6I4529_$1I4488_$1I4620_ADDRA[4], _6I4529_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_491_3 (_6I4529_$1I4488_$1I4620_ADDRA[3], _6I4529_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_491_2 (_6I4529_$1I4488_$1I4620_ADDRA[2], _6I4529_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_491_1 (_6I4529_$1I4488_$1I4620_ADDRA[1], _6I4529_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_491_0 (_6I4529_$1I4488_$1I4620_ADDRA[0], _6I4529_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _6I4529_$1I4488_$1I4620_ADDRB;
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_492_9 (_6I4529_$1I4488_$1I4620_ADDRB[9], _6I4529_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_492_8 (_6I4529_$1I4488_$1I4620_ADDRB[8], _6I4529_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_492_7 (_6I4529_$1I4488_$1I4620_ADDRB[7], _6I4529_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_492_6 (_6I4529_$1I4488_$1I4620_ADDRB[6], _6I4529_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_492_5 (_6I4529_$1I4488_$1I4620_ADDRB[5], _6I4529_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_492_4 (_6I4529_$1I4488_$1I4620_ADDRB[4], _6I4529_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_492_3 (_6I4529_$1I4488_$1I4620_ADDRB[3], _6I4529_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_492_2 (_6I4529_$1I4488_$1I4620_ADDRB[2], _6I4529_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_492_1 (_6I4529_$1I4488_$1I4620_ADDRB[1], _6I4529_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_492_0 (_6I4529_$1I4488_$1I4620_ADDRB[0], _6I4529_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _6I4529_$1I4488_$1I4620_CLKA;
 reg [1:16] _6I4529_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_493 (_6I4529_$1I4488_$1I4620_CLKA, _6I4529_$1I4488_$1I4620_CLKA__vlIN);

 wire  _6I4529_$1I4488_$1I4620_CLKB;
 reg [1:16] _6I4529_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_494 (_6I4529_$1I4488_$1I4620_CLKB, _6I4529_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _6I4529_$1I4488_$1I4620_DIA;
 reg [1:16] _6I4529_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_495_7 (_6I4529_$1I4488_$1I4620_DIA[7], _6I4529_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_495_6 (_6I4529_$1I4488_$1I4620_DIA[6], _6I4529_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_495_5 (_6I4529_$1I4488_$1I4620_DIA[5], _6I4529_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_495_4 (_6I4529_$1I4488_$1I4620_DIA[4], _6I4529_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_495_3 (_6I4529_$1I4488_$1I4620_DIA[3], _6I4529_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_495_2 (_6I4529_$1I4488_$1I4620_DIA[2], _6I4529_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_495_1 (_6I4529_$1I4488_$1I4620_DIA[1], _6I4529_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_495_0 (_6I4529_$1I4488_$1I4620_DIA[0], _6I4529_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _6I4529_$1I4488_$1I4620_DIB;
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_496_15 (_6I4529_$1I4488_$1I4620_DIB[15], _6I4529_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_496_14 (_6I4529_$1I4488_$1I4620_DIB[14], _6I4529_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_496_13 (_6I4529_$1I4488_$1I4620_DIB[13], _6I4529_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_496_12 (_6I4529_$1I4488_$1I4620_DIB[12], _6I4529_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_496_11 (_6I4529_$1I4488_$1I4620_DIB[11], _6I4529_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_496_10 (_6I4529_$1I4488_$1I4620_DIB[10], _6I4529_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_496_9 (_6I4529_$1I4488_$1I4620_DIB[9], _6I4529_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_496_8 (_6I4529_$1I4488_$1I4620_DIB[8], _6I4529_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_496_7 (_6I4529_$1I4488_$1I4620_DIB[7], _6I4529_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_496_6 (_6I4529_$1I4488_$1I4620_DIB[6], _6I4529_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_496_5 (_6I4529_$1I4488_$1I4620_DIB[5], _6I4529_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_496_4 (_6I4529_$1I4488_$1I4620_DIB[4], _6I4529_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_496_3 (_6I4529_$1I4488_$1I4620_DIB[3], _6I4529_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_496_2 (_6I4529_$1I4488_$1I4620_DIB[2], _6I4529_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_496_1 (_6I4529_$1I4488_$1I4620_DIB[1], _6I4529_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_496_0 (_6I4529_$1I4488_$1I4620_DIB[0], _6I4529_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _6I4529_$1I4488_$1I4620_DIPA;
 reg [1:16] _6I4529_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_497_0 (_6I4529_$1I4488_$1I4620_DIPA[0], _6I4529_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _6I4529_$1I4488_$1I4620_DIPB;
 reg [1:16] _6I4529_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_498_1 (_6I4529_$1I4488_$1I4620_DIPB[1], _6I4529_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _6I4529_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_498_0 (_6I4529_$1I4488_$1I4620_DIPB[0], _6I4529_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _6I4529_$1I4488_$1I4620_ENA;
 reg [1:16] _6I4529_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_499 (_6I4529_$1I4488_$1I4620_ENA, _6I4529_$1I4488_$1I4620_ENA__vlIN);

 wire  _6I4529_$1I4488_$1I4620_ENB;
 reg [1:16] _6I4529_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_500 (_6I4529_$1I4488_$1I4620_ENB, _6I4529_$1I4488_$1I4620_ENB__vlIN);

 wire  _6I4529_$1I4488_$1I4620_SSRA;
 reg [1:16] _6I4529_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_501 (_6I4529_$1I4488_$1I4620_SSRA, _6I4529_$1I4488_$1I4620_SSRA__vlIN);

 wire  _6I4529_$1I4488_$1I4620_SSRB;
 reg [1:16] _6I4529_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_502 (_6I4529_$1I4488_$1I4620_SSRB, _6I4529_$1I4488_$1I4620_SSRB__vlIN);

 wire  _6I4529_$1I4488_$1I4620_WEA;
 reg [1:16] _6I4529_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_503 (_6I4529_$1I4488_$1I4620_WEA, _6I4529_$1I4488_$1I4620_WEA__vlIN);

 wire  _6I4529_$1I4488_$1I4620_WEB;
 reg [1:16] _6I4529_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_504 (_6I4529_$1I4488_$1I4620_WEB, _6I4529_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _6I4529_$1I4488_$1I4620 ( _6I4529_$1I4488_$1I4620_DOA , _6I4529_$1I4488_$1I4620_DOB , _6I4529_$1I4488_$1I4620_DOPA , _6I4529_$1I4488_$1I4620_DOPB , _6I4529_$1I4488_$1I4620_ADDRA , _6I4529_$1I4488_$1I4620_ADDRB , _6I4529_$1I4488_$1I4620_CLKA , _6I4529_$1I4488_$1I4620_CLKB , _6I4529_$1I4488_$1I4620_DIA , _6I4529_$1I4488_$1I4620_DIB , _6I4529_$1I4488_$1I4620_DIPA , _6I4529_$1I4488_$1I4620_DIPB , _6I4529_$1I4488_$1I4620_ENA , _6I4529_$1I4488_$1I4620_ENB , _6I4529_$1I4488_$1I4620_SSRA , _6I4529_$1I4488_$1I4620_SSRB , _6I4529_$1I4488_$1I4620_WEA , _6I4529_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4504_$1I4488_$1I4621_DOA;

 wire [15:0] _6I4504_$1I4488_$1I4621_DOB;

 wire [0:0] _6I4504_$1I4488_$1I4621_DOPA;

 wire [1:0] _6I4504_$1I4488_$1I4621_DOPB;

 wire [10:0] _6I4504_$1I4488_$1I4621_ADDRA;
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_505_10 (_6I4504_$1I4488_$1I4621_ADDRA[10], _6I4504_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_505_9 (_6I4504_$1I4488_$1I4621_ADDRA[9], _6I4504_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_505_8 (_6I4504_$1I4488_$1I4621_ADDRA[8], _6I4504_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_505_7 (_6I4504_$1I4488_$1I4621_ADDRA[7], _6I4504_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_505_6 (_6I4504_$1I4488_$1I4621_ADDRA[6], _6I4504_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_505_5 (_6I4504_$1I4488_$1I4621_ADDRA[5], _6I4504_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_505_4 (_6I4504_$1I4488_$1I4621_ADDRA[4], _6I4504_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_505_3 (_6I4504_$1I4488_$1I4621_ADDRA[3], _6I4504_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_505_2 (_6I4504_$1I4488_$1I4621_ADDRA[2], _6I4504_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_505_1 (_6I4504_$1I4488_$1I4621_ADDRA[1], _6I4504_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_505_0 (_6I4504_$1I4488_$1I4621_ADDRA[0], _6I4504_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _6I4504_$1I4488_$1I4621_ADDRB;
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_506_9 (_6I4504_$1I4488_$1I4621_ADDRB[9], _6I4504_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_506_8 (_6I4504_$1I4488_$1I4621_ADDRB[8], _6I4504_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_506_7 (_6I4504_$1I4488_$1I4621_ADDRB[7], _6I4504_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_506_6 (_6I4504_$1I4488_$1I4621_ADDRB[6], _6I4504_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_506_5 (_6I4504_$1I4488_$1I4621_ADDRB[5], _6I4504_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_506_4 (_6I4504_$1I4488_$1I4621_ADDRB[4], _6I4504_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_506_3 (_6I4504_$1I4488_$1I4621_ADDRB[3], _6I4504_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_506_2 (_6I4504_$1I4488_$1I4621_ADDRB[2], _6I4504_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_506_1 (_6I4504_$1I4488_$1I4621_ADDRB[1], _6I4504_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_506_0 (_6I4504_$1I4488_$1I4621_ADDRB[0], _6I4504_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _6I4504_$1I4488_$1I4621_CLKA;
 reg [1:16] _6I4504_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_507 (_6I4504_$1I4488_$1I4621_CLKA, _6I4504_$1I4488_$1I4621_CLKA__vlIN);

 wire  _6I4504_$1I4488_$1I4621_CLKB;
 reg [1:16] _6I4504_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_508 (_6I4504_$1I4488_$1I4621_CLKB, _6I4504_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _6I4504_$1I4488_$1I4621_DIA;
 reg [1:16] _6I4504_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_509_7 (_6I4504_$1I4488_$1I4621_DIA[7], _6I4504_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_509_6 (_6I4504_$1I4488_$1I4621_DIA[6], _6I4504_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_509_5 (_6I4504_$1I4488_$1I4621_DIA[5], _6I4504_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_509_4 (_6I4504_$1I4488_$1I4621_DIA[4], _6I4504_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_509_3 (_6I4504_$1I4488_$1I4621_DIA[3], _6I4504_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_509_2 (_6I4504_$1I4488_$1I4621_DIA[2], _6I4504_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_509_1 (_6I4504_$1I4488_$1I4621_DIA[1], _6I4504_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_509_0 (_6I4504_$1I4488_$1I4621_DIA[0], _6I4504_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _6I4504_$1I4488_$1I4621_DIB;
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_510_15 (_6I4504_$1I4488_$1I4621_DIB[15], _6I4504_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_510_14 (_6I4504_$1I4488_$1I4621_DIB[14], _6I4504_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_510_13 (_6I4504_$1I4488_$1I4621_DIB[13], _6I4504_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_510_12 (_6I4504_$1I4488_$1I4621_DIB[12], _6I4504_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_510_11 (_6I4504_$1I4488_$1I4621_DIB[11], _6I4504_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_510_10 (_6I4504_$1I4488_$1I4621_DIB[10], _6I4504_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_510_9 (_6I4504_$1I4488_$1I4621_DIB[9], _6I4504_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_510_8 (_6I4504_$1I4488_$1I4621_DIB[8], _6I4504_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_510_7 (_6I4504_$1I4488_$1I4621_DIB[7], _6I4504_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_510_6 (_6I4504_$1I4488_$1I4621_DIB[6], _6I4504_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_510_5 (_6I4504_$1I4488_$1I4621_DIB[5], _6I4504_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_510_4 (_6I4504_$1I4488_$1I4621_DIB[4], _6I4504_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_510_3 (_6I4504_$1I4488_$1I4621_DIB[3], _6I4504_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_510_2 (_6I4504_$1I4488_$1I4621_DIB[2], _6I4504_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_510_1 (_6I4504_$1I4488_$1I4621_DIB[1], _6I4504_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_510_0 (_6I4504_$1I4488_$1I4621_DIB[0], _6I4504_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _6I4504_$1I4488_$1I4621_DIPA;
 reg [1:16] _6I4504_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_511_0 (_6I4504_$1I4488_$1I4621_DIPA[0], _6I4504_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _6I4504_$1I4488_$1I4621_DIPB;
 reg [1:16] _6I4504_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_512_1 (_6I4504_$1I4488_$1I4621_DIPB[1], _6I4504_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_512_0 (_6I4504_$1I4488_$1I4621_DIPB[0], _6I4504_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _6I4504_$1I4488_$1I4621_ENA;
 reg [1:16] _6I4504_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_513 (_6I4504_$1I4488_$1I4621_ENA, _6I4504_$1I4488_$1I4621_ENA__vlIN);

 wire  _6I4504_$1I4488_$1I4621_ENB;
 reg [1:16] _6I4504_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_514 (_6I4504_$1I4488_$1I4621_ENB, _6I4504_$1I4488_$1I4621_ENB__vlIN);

 wire  _6I4504_$1I4488_$1I4621_SSRA;
 reg [1:16] _6I4504_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_515 (_6I4504_$1I4488_$1I4621_SSRA, _6I4504_$1I4488_$1I4621_SSRA__vlIN);

 wire  _6I4504_$1I4488_$1I4621_SSRB;
 reg [1:16] _6I4504_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_516 (_6I4504_$1I4488_$1I4621_SSRB, _6I4504_$1I4488_$1I4621_SSRB__vlIN);

 wire  _6I4504_$1I4488_$1I4621_WEA;
 reg [1:16] _6I4504_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_517 (_6I4504_$1I4488_$1I4621_WEA, _6I4504_$1I4488_$1I4621_WEA__vlIN);

 wire  _6I4504_$1I4488_$1I4621_WEB;
 reg [1:16] _6I4504_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_518 (_6I4504_$1I4488_$1I4621_WEB, _6I4504_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _6I4504_$1I4488_$1I4621 ( _6I4504_$1I4488_$1I4621_DOA , _6I4504_$1I4488_$1I4621_DOB , _6I4504_$1I4488_$1I4621_DOPA , _6I4504_$1I4488_$1I4621_DOPB , _6I4504_$1I4488_$1I4621_ADDRA , _6I4504_$1I4488_$1I4621_ADDRB , _6I4504_$1I4488_$1I4621_CLKA , _6I4504_$1I4488_$1I4621_CLKB , _6I4504_$1I4488_$1I4621_DIA , _6I4504_$1I4488_$1I4621_DIB , _6I4504_$1I4488_$1I4621_DIPA , _6I4504_$1I4488_$1I4621_DIPB , _6I4504_$1I4488_$1I4621_ENA , _6I4504_$1I4488_$1I4621_ENB , _6I4504_$1I4488_$1I4621_SSRA , _6I4504_$1I4488_$1I4621_SSRB , _6I4504_$1I4488_$1I4621_WEA , _6I4504_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4504_$1I4488_$1I4620_DOA;

 wire [15:0] _6I4504_$1I4488_$1I4620_DOB;

 wire [0:0] _6I4504_$1I4488_$1I4620_DOPA;

 wire [1:0] _6I4504_$1I4488_$1I4620_DOPB;

 wire [10:0] _6I4504_$1I4488_$1I4620_ADDRA;
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_519_10 (_6I4504_$1I4488_$1I4620_ADDRA[10], _6I4504_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_519_9 (_6I4504_$1I4488_$1I4620_ADDRA[9], _6I4504_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_519_8 (_6I4504_$1I4488_$1I4620_ADDRA[8], _6I4504_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_519_7 (_6I4504_$1I4488_$1I4620_ADDRA[7], _6I4504_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_519_6 (_6I4504_$1I4488_$1I4620_ADDRA[6], _6I4504_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_519_5 (_6I4504_$1I4488_$1I4620_ADDRA[5], _6I4504_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_519_4 (_6I4504_$1I4488_$1I4620_ADDRA[4], _6I4504_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_519_3 (_6I4504_$1I4488_$1I4620_ADDRA[3], _6I4504_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_519_2 (_6I4504_$1I4488_$1I4620_ADDRA[2], _6I4504_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_519_1 (_6I4504_$1I4488_$1I4620_ADDRA[1], _6I4504_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_519_0 (_6I4504_$1I4488_$1I4620_ADDRA[0], _6I4504_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _6I4504_$1I4488_$1I4620_ADDRB;
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_520_9 (_6I4504_$1I4488_$1I4620_ADDRB[9], _6I4504_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_520_8 (_6I4504_$1I4488_$1I4620_ADDRB[8], _6I4504_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_520_7 (_6I4504_$1I4488_$1I4620_ADDRB[7], _6I4504_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_520_6 (_6I4504_$1I4488_$1I4620_ADDRB[6], _6I4504_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_520_5 (_6I4504_$1I4488_$1I4620_ADDRB[5], _6I4504_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_520_4 (_6I4504_$1I4488_$1I4620_ADDRB[4], _6I4504_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_520_3 (_6I4504_$1I4488_$1I4620_ADDRB[3], _6I4504_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_520_2 (_6I4504_$1I4488_$1I4620_ADDRB[2], _6I4504_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_520_1 (_6I4504_$1I4488_$1I4620_ADDRB[1], _6I4504_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_520_0 (_6I4504_$1I4488_$1I4620_ADDRB[0], _6I4504_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _6I4504_$1I4488_$1I4620_CLKA;
 reg [1:16] _6I4504_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_521 (_6I4504_$1I4488_$1I4620_CLKA, _6I4504_$1I4488_$1I4620_CLKA__vlIN);

 wire  _6I4504_$1I4488_$1I4620_CLKB;
 reg [1:16] _6I4504_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_522 (_6I4504_$1I4488_$1I4620_CLKB, _6I4504_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _6I4504_$1I4488_$1I4620_DIA;
 reg [1:16] _6I4504_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_523_7 (_6I4504_$1I4488_$1I4620_DIA[7], _6I4504_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_523_6 (_6I4504_$1I4488_$1I4620_DIA[6], _6I4504_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_523_5 (_6I4504_$1I4488_$1I4620_DIA[5], _6I4504_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_523_4 (_6I4504_$1I4488_$1I4620_DIA[4], _6I4504_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_523_3 (_6I4504_$1I4488_$1I4620_DIA[3], _6I4504_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_523_2 (_6I4504_$1I4488_$1I4620_DIA[2], _6I4504_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_523_1 (_6I4504_$1I4488_$1I4620_DIA[1], _6I4504_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_523_0 (_6I4504_$1I4488_$1I4620_DIA[0], _6I4504_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _6I4504_$1I4488_$1I4620_DIB;
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_524_15 (_6I4504_$1I4488_$1I4620_DIB[15], _6I4504_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_524_14 (_6I4504_$1I4488_$1I4620_DIB[14], _6I4504_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_524_13 (_6I4504_$1I4488_$1I4620_DIB[13], _6I4504_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_524_12 (_6I4504_$1I4488_$1I4620_DIB[12], _6I4504_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_524_11 (_6I4504_$1I4488_$1I4620_DIB[11], _6I4504_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_524_10 (_6I4504_$1I4488_$1I4620_DIB[10], _6I4504_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_524_9 (_6I4504_$1I4488_$1I4620_DIB[9], _6I4504_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_524_8 (_6I4504_$1I4488_$1I4620_DIB[8], _6I4504_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_524_7 (_6I4504_$1I4488_$1I4620_DIB[7], _6I4504_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_524_6 (_6I4504_$1I4488_$1I4620_DIB[6], _6I4504_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_524_5 (_6I4504_$1I4488_$1I4620_DIB[5], _6I4504_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_524_4 (_6I4504_$1I4488_$1I4620_DIB[4], _6I4504_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_524_3 (_6I4504_$1I4488_$1I4620_DIB[3], _6I4504_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_524_2 (_6I4504_$1I4488_$1I4620_DIB[2], _6I4504_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_524_1 (_6I4504_$1I4488_$1I4620_DIB[1], _6I4504_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_524_0 (_6I4504_$1I4488_$1I4620_DIB[0], _6I4504_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _6I4504_$1I4488_$1I4620_DIPA;
 reg [1:16] _6I4504_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_525_0 (_6I4504_$1I4488_$1I4620_DIPA[0], _6I4504_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _6I4504_$1I4488_$1I4620_DIPB;
 reg [1:16] _6I4504_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_526_1 (_6I4504_$1I4488_$1I4620_DIPB[1], _6I4504_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _6I4504_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_526_0 (_6I4504_$1I4488_$1I4620_DIPB[0], _6I4504_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _6I4504_$1I4488_$1I4620_ENA;
 reg [1:16] _6I4504_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_527 (_6I4504_$1I4488_$1I4620_ENA, _6I4504_$1I4488_$1I4620_ENA__vlIN);

 wire  _6I4504_$1I4488_$1I4620_ENB;
 reg [1:16] _6I4504_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_528 (_6I4504_$1I4488_$1I4620_ENB, _6I4504_$1I4488_$1I4620_ENB__vlIN);

 wire  _6I4504_$1I4488_$1I4620_SSRA;
 reg [1:16] _6I4504_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_529 (_6I4504_$1I4488_$1I4620_SSRA, _6I4504_$1I4488_$1I4620_SSRA__vlIN);

 wire  _6I4504_$1I4488_$1I4620_SSRB;
 reg [1:16] _6I4504_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_530 (_6I4504_$1I4488_$1I4620_SSRB, _6I4504_$1I4488_$1I4620_SSRB__vlIN);

 wire  _6I4504_$1I4488_$1I4620_WEA;
 reg [1:16] _6I4504_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_531 (_6I4504_$1I4488_$1I4620_WEA, _6I4504_$1I4488_$1I4620_WEA__vlIN);

 wire  _6I4504_$1I4488_$1I4620_WEB;
 reg [1:16] _6I4504_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_532 (_6I4504_$1I4488_$1I4620_WEB, _6I4504_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _6I4504_$1I4488_$1I4620 ( _6I4504_$1I4488_$1I4620_DOA , _6I4504_$1I4488_$1I4620_DOB , _6I4504_$1I4488_$1I4620_DOPA , _6I4504_$1I4488_$1I4620_DOPB , _6I4504_$1I4488_$1I4620_ADDRA , _6I4504_$1I4488_$1I4620_ADDRB , _6I4504_$1I4488_$1I4620_CLKA , _6I4504_$1I4488_$1I4620_CLKB , _6I4504_$1I4488_$1I4620_DIA , _6I4504_$1I4488_$1I4620_DIB , _6I4504_$1I4488_$1I4620_DIPA , _6I4504_$1I4488_$1I4620_DIPB , _6I4504_$1I4488_$1I4620_ENA , _6I4504_$1I4488_$1I4620_ENB , _6I4504_$1I4488_$1I4620_SSRA , _6I4504_$1I4488_$1I4620_SSRB , _6I4504_$1I4488_$1I4620_WEA , _6I4504_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4479_$1I4488_$1I4621_DOA;

 wire [15:0] _6I4479_$1I4488_$1I4621_DOB;

 wire [0:0] _6I4479_$1I4488_$1I4621_DOPA;

 wire [1:0] _6I4479_$1I4488_$1I4621_DOPB;

 wire [10:0] _6I4479_$1I4488_$1I4621_ADDRA;
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_533_10 (_6I4479_$1I4488_$1I4621_ADDRA[10], _6I4479_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_533_9 (_6I4479_$1I4488_$1I4621_ADDRA[9], _6I4479_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_533_8 (_6I4479_$1I4488_$1I4621_ADDRA[8], _6I4479_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_533_7 (_6I4479_$1I4488_$1I4621_ADDRA[7], _6I4479_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_533_6 (_6I4479_$1I4488_$1I4621_ADDRA[6], _6I4479_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_533_5 (_6I4479_$1I4488_$1I4621_ADDRA[5], _6I4479_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_533_4 (_6I4479_$1I4488_$1I4621_ADDRA[4], _6I4479_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_533_3 (_6I4479_$1I4488_$1I4621_ADDRA[3], _6I4479_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_533_2 (_6I4479_$1I4488_$1I4621_ADDRA[2], _6I4479_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_533_1 (_6I4479_$1I4488_$1I4621_ADDRA[1], _6I4479_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_533_0 (_6I4479_$1I4488_$1I4621_ADDRA[0], _6I4479_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _6I4479_$1I4488_$1I4621_ADDRB;
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_534_9 (_6I4479_$1I4488_$1I4621_ADDRB[9], _6I4479_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_534_8 (_6I4479_$1I4488_$1I4621_ADDRB[8], _6I4479_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_534_7 (_6I4479_$1I4488_$1I4621_ADDRB[7], _6I4479_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_534_6 (_6I4479_$1I4488_$1I4621_ADDRB[6], _6I4479_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_534_5 (_6I4479_$1I4488_$1I4621_ADDRB[5], _6I4479_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_534_4 (_6I4479_$1I4488_$1I4621_ADDRB[4], _6I4479_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_534_3 (_6I4479_$1I4488_$1I4621_ADDRB[3], _6I4479_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_534_2 (_6I4479_$1I4488_$1I4621_ADDRB[2], _6I4479_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_534_1 (_6I4479_$1I4488_$1I4621_ADDRB[1], _6I4479_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_534_0 (_6I4479_$1I4488_$1I4621_ADDRB[0], _6I4479_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _6I4479_$1I4488_$1I4621_CLKA;
 reg [1:16] _6I4479_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_535 (_6I4479_$1I4488_$1I4621_CLKA, _6I4479_$1I4488_$1I4621_CLKA__vlIN);

 wire  _6I4479_$1I4488_$1I4621_CLKB;
 reg [1:16] _6I4479_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_536 (_6I4479_$1I4488_$1I4621_CLKB, _6I4479_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _6I4479_$1I4488_$1I4621_DIA;
 reg [1:16] _6I4479_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_537_7 (_6I4479_$1I4488_$1I4621_DIA[7], _6I4479_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_537_6 (_6I4479_$1I4488_$1I4621_DIA[6], _6I4479_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_537_5 (_6I4479_$1I4488_$1I4621_DIA[5], _6I4479_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_537_4 (_6I4479_$1I4488_$1I4621_DIA[4], _6I4479_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_537_3 (_6I4479_$1I4488_$1I4621_DIA[3], _6I4479_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_537_2 (_6I4479_$1I4488_$1I4621_DIA[2], _6I4479_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_537_1 (_6I4479_$1I4488_$1I4621_DIA[1], _6I4479_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_537_0 (_6I4479_$1I4488_$1I4621_DIA[0], _6I4479_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _6I4479_$1I4488_$1I4621_DIB;
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_538_15 (_6I4479_$1I4488_$1I4621_DIB[15], _6I4479_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_538_14 (_6I4479_$1I4488_$1I4621_DIB[14], _6I4479_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_538_13 (_6I4479_$1I4488_$1I4621_DIB[13], _6I4479_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_538_12 (_6I4479_$1I4488_$1I4621_DIB[12], _6I4479_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_538_11 (_6I4479_$1I4488_$1I4621_DIB[11], _6I4479_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_538_10 (_6I4479_$1I4488_$1I4621_DIB[10], _6I4479_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_538_9 (_6I4479_$1I4488_$1I4621_DIB[9], _6I4479_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_538_8 (_6I4479_$1I4488_$1I4621_DIB[8], _6I4479_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_538_7 (_6I4479_$1I4488_$1I4621_DIB[7], _6I4479_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_538_6 (_6I4479_$1I4488_$1I4621_DIB[6], _6I4479_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_538_5 (_6I4479_$1I4488_$1I4621_DIB[5], _6I4479_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_538_4 (_6I4479_$1I4488_$1I4621_DIB[4], _6I4479_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_538_3 (_6I4479_$1I4488_$1I4621_DIB[3], _6I4479_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_538_2 (_6I4479_$1I4488_$1I4621_DIB[2], _6I4479_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_538_1 (_6I4479_$1I4488_$1I4621_DIB[1], _6I4479_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_538_0 (_6I4479_$1I4488_$1I4621_DIB[0], _6I4479_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _6I4479_$1I4488_$1I4621_DIPA;
 reg [1:16] _6I4479_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_539_0 (_6I4479_$1I4488_$1I4621_DIPA[0], _6I4479_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _6I4479_$1I4488_$1I4621_DIPB;
 reg [1:16] _6I4479_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_540_1 (_6I4479_$1I4488_$1I4621_DIPB[1], _6I4479_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_540_0 (_6I4479_$1I4488_$1I4621_DIPB[0], _6I4479_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _6I4479_$1I4488_$1I4621_ENA;
 reg [1:16] _6I4479_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_541 (_6I4479_$1I4488_$1I4621_ENA, _6I4479_$1I4488_$1I4621_ENA__vlIN);

 wire  _6I4479_$1I4488_$1I4621_ENB;
 reg [1:16] _6I4479_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_542 (_6I4479_$1I4488_$1I4621_ENB, _6I4479_$1I4488_$1I4621_ENB__vlIN);

 wire  _6I4479_$1I4488_$1I4621_SSRA;
 reg [1:16] _6I4479_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_543 (_6I4479_$1I4488_$1I4621_SSRA, _6I4479_$1I4488_$1I4621_SSRA__vlIN);

 wire  _6I4479_$1I4488_$1I4621_SSRB;
 reg [1:16] _6I4479_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_544 (_6I4479_$1I4488_$1I4621_SSRB, _6I4479_$1I4488_$1I4621_SSRB__vlIN);

 wire  _6I4479_$1I4488_$1I4621_WEA;
 reg [1:16] _6I4479_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_545 (_6I4479_$1I4488_$1I4621_WEA, _6I4479_$1I4488_$1I4621_WEA__vlIN);

 wire  _6I4479_$1I4488_$1I4621_WEB;
 reg [1:16] _6I4479_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_546 (_6I4479_$1I4488_$1I4621_WEB, _6I4479_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _6I4479_$1I4488_$1I4621 ( _6I4479_$1I4488_$1I4621_DOA , _6I4479_$1I4488_$1I4621_DOB , _6I4479_$1I4488_$1I4621_DOPA , _6I4479_$1I4488_$1I4621_DOPB , _6I4479_$1I4488_$1I4621_ADDRA , _6I4479_$1I4488_$1I4621_ADDRB , _6I4479_$1I4488_$1I4621_CLKA , _6I4479_$1I4488_$1I4621_CLKB , _6I4479_$1I4488_$1I4621_DIA , _6I4479_$1I4488_$1I4621_DIB , _6I4479_$1I4488_$1I4621_DIPA , _6I4479_$1I4488_$1I4621_DIPB , _6I4479_$1I4488_$1I4621_ENA , _6I4479_$1I4488_$1I4621_ENB , _6I4479_$1I4488_$1I4621_SSRA , _6I4479_$1I4488_$1I4621_SSRB , _6I4479_$1I4488_$1I4621_WEA , _6I4479_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4479_$1I4488_$1I4620_DOA;

 wire [15:0] _6I4479_$1I4488_$1I4620_DOB;

 wire [0:0] _6I4479_$1I4488_$1I4620_DOPA;

 wire [1:0] _6I4479_$1I4488_$1I4620_DOPB;

 wire [10:0] _6I4479_$1I4488_$1I4620_ADDRA;
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_547_10 (_6I4479_$1I4488_$1I4620_ADDRA[10], _6I4479_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_547_9 (_6I4479_$1I4488_$1I4620_ADDRA[9], _6I4479_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_547_8 (_6I4479_$1I4488_$1I4620_ADDRA[8], _6I4479_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_547_7 (_6I4479_$1I4488_$1I4620_ADDRA[7], _6I4479_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_547_6 (_6I4479_$1I4488_$1I4620_ADDRA[6], _6I4479_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_547_5 (_6I4479_$1I4488_$1I4620_ADDRA[5], _6I4479_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_547_4 (_6I4479_$1I4488_$1I4620_ADDRA[4], _6I4479_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_547_3 (_6I4479_$1I4488_$1I4620_ADDRA[3], _6I4479_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_547_2 (_6I4479_$1I4488_$1I4620_ADDRA[2], _6I4479_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_547_1 (_6I4479_$1I4488_$1I4620_ADDRA[1], _6I4479_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_547_0 (_6I4479_$1I4488_$1I4620_ADDRA[0], _6I4479_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _6I4479_$1I4488_$1I4620_ADDRB;
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_548_9 (_6I4479_$1I4488_$1I4620_ADDRB[9], _6I4479_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_548_8 (_6I4479_$1I4488_$1I4620_ADDRB[8], _6I4479_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_548_7 (_6I4479_$1I4488_$1I4620_ADDRB[7], _6I4479_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_548_6 (_6I4479_$1I4488_$1I4620_ADDRB[6], _6I4479_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_548_5 (_6I4479_$1I4488_$1I4620_ADDRB[5], _6I4479_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_548_4 (_6I4479_$1I4488_$1I4620_ADDRB[4], _6I4479_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_548_3 (_6I4479_$1I4488_$1I4620_ADDRB[3], _6I4479_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_548_2 (_6I4479_$1I4488_$1I4620_ADDRB[2], _6I4479_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_548_1 (_6I4479_$1I4488_$1I4620_ADDRB[1], _6I4479_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_548_0 (_6I4479_$1I4488_$1I4620_ADDRB[0], _6I4479_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _6I4479_$1I4488_$1I4620_CLKA;
 reg [1:16] _6I4479_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_549 (_6I4479_$1I4488_$1I4620_CLKA, _6I4479_$1I4488_$1I4620_CLKA__vlIN);

 wire  _6I4479_$1I4488_$1I4620_CLKB;
 reg [1:16] _6I4479_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_550 (_6I4479_$1I4488_$1I4620_CLKB, _6I4479_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _6I4479_$1I4488_$1I4620_DIA;
 reg [1:16] _6I4479_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_551_7 (_6I4479_$1I4488_$1I4620_DIA[7], _6I4479_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_551_6 (_6I4479_$1I4488_$1I4620_DIA[6], _6I4479_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_551_5 (_6I4479_$1I4488_$1I4620_DIA[5], _6I4479_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_551_4 (_6I4479_$1I4488_$1I4620_DIA[4], _6I4479_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_551_3 (_6I4479_$1I4488_$1I4620_DIA[3], _6I4479_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_551_2 (_6I4479_$1I4488_$1I4620_DIA[2], _6I4479_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_551_1 (_6I4479_$1I4488_$1I4620_DIA[1], _6I4479_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_551_0 (_6I4479_$1I4488_$1I4620_DIA[0], _6I4479_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _6I4479_$1I4488_$1I4620_DIB;
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_552_15 (_6I4479_$1I4488_$1I4620_DIB[15], _6I4479_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_552_14 (_6I4479_$1I4488_$1I4620_DIB[14], _6I4479_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_552_13 (_6I4479_$1I4488_$1I4620_DIB[13], _6I4479_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_552_12 (_6I4479_$1I4488_$1I4620_DIB[12], _6I4479_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_552_11 (_6I4479_$1I4488_$1I4620_DIB[11], _6I4479_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_552_10 (_6I4479_$1I4488_$1I4620_DIB[10], _6I4479_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_552_9 (_6I4479_$1I4488_$1I4620_DIB[9], _6I4479_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_552_8 (_6I4479_$1I4488_$1I4620_DIB[8], _6I4479_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_552_7 (_6I4479_$1I4488_$1I4620_DIB[7], _6I4479_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_552_6 (_6I4479_$1I4488_$1I4620_DIB[6], _6I4479_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_552_5 (_6I4479_$1I4488_$1I4620_DIB[5], _6I4479_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_552_4 (_6I4479_$1I4488_$1I4620_DIB[4], _6I4479_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_552_3 (_6I4479_$1I4488_$1I4620_DIB[3], _6I4479_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_552_2 (_6I4479_$1I4488_$1I4620_DIB[2], _6I4479_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_552_1 (_6I4479_$1I4488_$1I4620_DIB[1], _6I4479_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_552_0 (_6I4479_$1I4488_$1I4620_DIB[0], _6I4479_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _6I4479_$1I4488_$1I4620_DIPA;
 reg [1:16] _6I4479_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_553_0 (_6I4479_$1I4488_$1I4620_DIPA[0], _6I4479_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _6I4479_$1I4488_$1I4620_DIPB;
 reg [1:16] _6I4479_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_554_1 (_6I4479_$1I4488_$1I4620_DIPB[1], _6I4479_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _6I4479_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_554_0 (_6I4479_$1I4488_$1I4620_DIPB[0], _6I4479_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _6I4479_$1I4488_$1I4620_ENA;
 reg [1:16] _6I4479_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_555 (_6I4479_$1I4488_$1I4620_ENA, _6I4479_$1I4488_$1I4620_ENA__vlIN);

 wire  _6I4479_$1I4488_$1I4620_ENB;
 reg [1:16] _6I4479_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_556 (_6I4479_$1I4488_$1I4620_ENB, _6I4479_$1I4488_$1I4620_ENB__vlIN);

 wire  _6I4479_$1I4488_$1I4620_SSRA;
 reg [1:16] _6I4479_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_557 (_6I4479_$1I4488_$1I4620_SSRA, _6I4479_$1I4488_$1I4620_SSRA__vlIN);

 wire  _6I4479_$1I4488_$1I4620_SSRB;
 reg [1:16] _6I4479_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_558 (_6I4479_$1I4488_$1I4620_SSRB, _6I4479_$1I4488_$1I4620_SSRB__vlIN);

 wire  _6I4479_$1I4488_$1I4620_WEA;
 reg [1:16] _6I4479_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_559 (_6I4479_$1I4488_$1I4620_WEA, _6I4479_$1I4488_$1I4620_WEA__vlIN);

 wire  _6I4479_$1I4488_$1I4620_WEB;
 reg [1:16] _6I4479_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_560 (_6I4479_$1I4488_$1I4620_WEB, _6I4479_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _6I4479_$1I4488_$1I4620 ( _6I4479_$1I4488_$1I4620_DOA , _6I4479_$1I4488_$1I4620_DOB , _6I4479_$1I4488_$1I4620_DOPA , _6I4479_$1I4488_$1I4620_DOPB , _6I4479_$1I4488_$1I4620_ADDRA , _6I4479_$1I4488_$1I4620_ADDRB , _6I4479_$1I4488_$1I4620_CLKA , _6I4479_$1I4488_$1I4620_CLKB , _6I4479_$1I4488_$1I4620_DIA , _6I4479_$1I4488_$1I4620_DIB , _6I4479_$1I4488_$1I4620_DIPA , _6I4479_$1I4488_$1I4620_DIPB , _6I4479_$1I4488_$1I4620_ENA , _6I4479_$1I4488_$1I4620_ENB , _6I4479_$1I4488_$1I4620_SSRA , _6I4479_$1I4488_$1I4620_SSRB , _6I4479_$1I4488_$1I4620_WEA , _6I4479_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [4:0] _6I4446_$1I4152_din;
 reg [1:16] _6I4446_$1I4152_din_4__vlIN;
 cstw cstw_561_4 (_6I4446_$1I4152_din[4], _6I4446_$1I4152_din_4__vlIN);
 reg [1:16] _6I4446_$1I4152_din_3__vlIN;
 cstw cstw_561_3 (_6I4446_$1I4152_din[3], _6I4446_$1I4152_din_3__vlIN);
 reg [1:16] _6I4446_$1I4152_din_2__vlIN;
 cstw cstw_561_2 (_6I4446_$1I4152_din[2], _6I4446_$1I4152_din_2__vlIN);
 reg [1:16] _6I4446_$1I4152_din_1__vlIN;
 cstw cstw_561_1 (_6I4446_$1I4152_din[1], _6I4446_$1I4152_din_1__vlIN);
 reg [1:16] _6I4446_$1I4152_din_0__vlIN;
 cstw cstw_561_0 (_6I4446_$1I4152_din[0], _6I4446_$1I4152_din_0__vlIN);

 wire  _6I4446_$1I4152_wr_en;
 reg [1:16] _6I4446_$1I4152_wr_en__vlIN;
 cstw cstw_562 (_6I4446_$1I4152_wr_en, _6I4446_$1I4152_wr_en__vlIN);

 wire  _6I4446_$1I4152_wr_clk;
 reg [1:16] _6I4446_$1I4152_wr_clk__vlIN;
 cstw cstw_563 (_6I4446_$1I4152_wr_clk, _6I4446_$1I4152_wr_clk__vlIN);

 wire  _6I4446_$1I4152_rd_en;
 reg [1:16] _6I4446_$1I4152_rd_en__vlIN;
 cstw cstw_564 (_6I4446_$1I4152_rd_en, _6I4446_$1I4152_rd_en__vlIN);

 wire  _6I4446_$1I4152_rd_clk;
 reg [1:16] _6I4446_$1I4152_rd_clk__vlIN;
 cstw cstw_565 (_6I4446_$1I4152_rd_clk, _6I4446_$1I4152_rd_clk__vlIN);

 wire  _6I4446_$1I4152_ainit;
 reg [1:16] _6I4446_$1I4152_ainit__vlIN;
 cstw cstw_566 (_6I4446_$1I4152_ainit, _6I4446_$1I4152_ainit__vlIN);

 wire [4:0] _6I4446_$1I4152_dout;

 wire  _6I4446_$1I4152_full;

 wire  _6I4446_$1I4152_empty;

 af_clb_5x31rpm _6I4446_$1I4152 ( _6I4446_$1I4152_din , _6I4446_$1I4152_wr_en , _6I4446_$1I4152_wr_clk , _6I4446_$1I4152_rd_en , _6I4446_$1I4152_rd_clk , _6I4446_$1I4152_ainit , _6I4446_$1I4152_dout , _6I4446_$1I4152_full , _6I4446_$1I4152_empty  );

// ----------------------------------- //

 wire  _6I4446_$1I3863_CHBONDDONE;

 wire [3:0] _6I4446_$1I3863_CHBONDO;

 wire  _6I4446_$1I3863_CONFIGOUT;

 wire [1:0] _6I4446_$1I3863_RXBUFSTATUS;

 wire [3:0] _6I4446_$1I3863_RXCHARISCOMMA;

 wire [3:0] _6I4446_$1I3863_RXCHARISK;

 wire  _6I4446_$1I3863_RXCHECKINGCRC;

 wire [2:0] _6I4446_$1I3863_RXCLKCORCNT;

 wire  _6I4446_$1I3863_RXCOMMADET;

 wire  _6I4446_$1I3863_RXCRCERR;

 wire [31:0] _6I4446_$1I3863_RXDATA;

 wire [3:0] _6I4446_$1I3863_RXDISPERR;

 wire [1:0] _6I4446_$1I3863_RXLOSSOFSYNC;

 wire [3:0] _6I4446_$1I3863_RXNOTINTABLE;

 wire  _6I4446_$1I3863_RXREALIGN;

 wire  _6I4446_$1I3863_RXRECCLK;

 wire [3:0] _6I4446_$1I3863_RXRUNDISP;

 wire  _6I4446_$1I3863_TXBUFERR;

 wire [3:0] _6I4446_$1I3863_TXKERR;

 wire  _6I4446_$1I3863_TXN;

 wire  _6I4446_$1I3863_TXP;

 wire [3:0] _6I4446_$1I3863_TXRUNDISP;

 wire  _6I4446_$1I3863_BREFCLK;
 reg [1:16] _6I4446_$1I3863_BREFCLK__vlIN;
 cstw cstw_567 (_6I4446_$1I3863_BREFCLK, _6I4446_$1I3863_BREFCLK__vlIN);

 wire  _6I4446_$1I3863_BREFCLK2;
 reg [1:16] _6I4446_$1I3863_BREFCLK2__vlIN;
 cstw cstw_568 (_6I4446_$1I3863_BREFCLK2, _6I4446_$1I3863_BREFCLK2__vlIN);

 wire [3:0] _6I4446_$1I3863_CHBONDI;
 reg [1:16] _6I4446_$1I3863_CHBONDI_3__vlIN;
 cstw cstw_569_3 (_6I4446_$1I3863_CHBONDI[3], _6I4446_$1I3863_CHBONDI_3__vlIN);
 reg [1:16] _6I4446_$1I3863_CHBONDI_2__vlIN;
 cstw cstw_569_2 (_6I4446_$1I3863_CHBONDI[2], _6I4446_$1I3863_CHBONDI_2__vlIN);
 reg [1:16] _6I4446_$1I3863_CHBONDI_1__vlIN;
 cstw cstw_569_1 (_6I4446_$1I3863_CHBONDI[1], _6I4446_$1I3863_CHBONDI_1__vlIN);
 reg [1:16] _6I4446_$1I3863_CHBONDI_0__vlIN;
 cstw cstw_569_0 (_6I4446_$1I3863_CHBONDI[0], _6I4446_$1I3863_CHBONDI_0__vlIN);

 wire  _6I4446_$1I3863_CONFIGENABLE;
 reg [1:16] _6I4446_$1I3863_CONFIGENABLE__vlIN;
 cstw cstw_570 (_6I4446_$1I3863_CONFIGENABLE, _6I4446_$1I3863_CONFIGENABLE__vlIN);

 wire  _6I4446_$1I3863_CONFIGIN;
 reg [1:16] _6I4446_$1I3863_CONFIGIN__vlIN;
 cstw cstw_571 (_6I4446_$1I3863_CONFIGIN, _6I4446_$1I3863_CONFIGIN__vlIN);

 wire  _6I4446_$1I3863_ENCHANSYNC;
 reg [1:16] _6I4446_$1I3863_ENCHANSYNC__vlIN;
 cstw cstw_572 (_6I4446_$1I3863_ENCHANSYNC, _6I4446_$1I3863_ENCHANSYNC__vlIN);

 wire  _6I4446_$1I3863_ENMCOMMAALIGN;
 reg [1:16] _6I4446_$1I3863_ENMCOMMAALIGN__vlIN;
 cstw cstw_573 (_6I4446_$1I3863_ENMCOMMAALIGN, _6I4446_$1I3863_ENMCOMMAALIGN__vlIN);

 wire  _6I4446_$1I3863_ENPCOMMAALIGN;
 reg [1:16] _6I4446_$1I3863_ENPCOMMAALIGN__vlIN;
 cstw cstw_574 (_6I4446_$1I3863_ENPCOMMAALIGN, _6I4446_$1I3863_ENPCOMMAALIGN__vlIN);

 wire [1:0] _6I4446_$1I3863_LOOPBACK;
 reg [1:16] _6I4446_$1I3863_LOOPBACK_1__vlIN;
 cstw cstw_575_1 (_6I4446_$1I3863_LOOPBACK[1], _6I4446_$1I3863_LOOPBACK_1__vlIN);
 reg [1:16] _6I4446_$1I3863_LOOPBACK_0__vlIN;
 cstw cstw_575_0 (_6I4446_$1I3863_LOOPBACK[0], _6I4446_$1I3863_LOOPBACK_0__vlIN);

 wire  _6I4446_$1I3863_POWERDOWN;
 reg [1:16] _6I4446_$1I3863_POWERDOWN__vlIN;
 cstw cstw_576 (_6I4446_$1I3863_POWERDOWN, _6I4446_$1I3863_POWERDOWN__vlIN);

 wire  _6I4446_$1I3863_REFCLK;
 reg [1:16] _6I4446_$1I3863_REFCLK__vlIN;
 cstw cstw_577 (_6I4446_$1I3863_REFCLK, _6I4446_$1I3863_REFCLK__vlIN);

 wire  _6I4446_$1I3863_REFCLK2;
 reg [1:16] _6I4446_$1I3863_REFCLK2__vlIN;
 cstw cstw_578 (_6I4446_$1I3863_REFCLK2, _6I4446_$1I3863_REFCLK2__vlIN);

 wire  _6I4446_$1I3863_REFCLKSEL;
 reg [1:16] _6I4446_$1I3863_REFCLKSEL__vlIN;
 cstw cstw_579 (_6I4446_$1I3863_REFCLKSEL, _6I4446_$1I3863_REFCLKSEL__vlIN);

 wire  _6I4446_$1I3863_RXN;
 reg [1:16] _6I4446_$1I3863_RXN__vlIN;
 cstw cstw_580 (_6I4446_$1I3863_RXN, _6I4446_$1I3863_RXN__vlIN);

 wire  _6I4446_$1I3863_RXP;
 reg [1:16] _6I4446_$1I3863_RXP__vlIN;
 cstw cstw_581 (_6I4446_$1I3863_RXP, _6I4446_$1I3863_RXP__vlIN);

 wire  _6I4446_$1I3863_RXPOLARITY;
 reg [1:16] _6I4446_$1I3863_RXPOLARITY__vlIN;
 cstw cstw_582 (_6I4446_$1I3863_RXPOLARITY, _6I4446_$1I3863_RXPOLARITY__vlIN);

 wire  _6I4446_$1I3863_RXRESET;
 reg [1:16] _6I4446_$1I3863_RXRESET__vlIN;
 cstw cstw_583 (_6I4446_$1I3863_RXRESET, _6I4446_$1I3863_RXRESET__vlIN);

 wire  _6I4446_$1I3863_RXUSRCLK;
 reg [1:16] _6I4446_$1I3863_RXUSRCLK__vlIN;
 cstw cstw_584 (_6I4446_$1I3863_RXUSRCLK, _6I4446_$1I3863_RXUSRCLK__vlIN);

 wire  _6I4446_$1I3863_RXUSRCLK2;
 reg [1:16] _6I4446_$1I3863_RXUSRCLK2__vlIN;
 cstw cstw_585 (_6I4446_$1I3863_RXUSRCLK2, _6I4446_$1I3863_RXUSRCLK2__vlIN);

 wire [3:0] _6I4446_$1I3863_TXBYPASS8B10B;
 reg [1:16] _6I4446_$1I3863_TXBYPASS8B10B_3__vlIN;
 cstw cstw_586_3 (_6I4446_$1I3863_TXBYPASS8B10B[3], _6I4446_$1I3863_TXBYPASS8B10B_3__vlIN);
 reg [1:16] _6I4446_$1I3863_TXBYPASS8B10B_2__vlIN;
 cstw cstw_586_2 (_6I4446_$1I3863_TXBYPASS8B10B[2], _6I4446_$1I3863_TXBYPASS8B10B_2__vlIN);
 reg [1:16] _6I4446_$1I3863_TXBYPASS8B10B_1__vlIN;
 cstw cstw_586_1 (_6I4446_$1I3863_TXBYPASS8B10B[1], _6I4446_$1I3863_TXBYPASS8B10B_1__vlIN);
 reg [1:16] _6I4446_$1I3863_TXBYPASS8B10B_0__vlIN;
 cstw cstw_586_0 (_6I4446_$1I3863_TXBYPASS8B10B[0], _6I4446_$1I3863_TXBYPASS8B10B_0__vlIN);

 wire [3:0] _6I4446_$1I3863_TXCHARDISPMODE;
 reg [1:16] _6I4446_$1I3863_TXCHARDISPMODE_3__vlIN;
 cstw cstw_587_3 (_6I4446_$1I3863_TXCHARDISPMODE[3], _6I4446_$1I3863_TXCHARDISPMODE_3__vlIN);
 reg [1:16] _6I4446_$1I3863_TXCHARDISPMODE_2__vlIN;
 cstw cstw_587_2 (_6I4446_$1I3863_TXCHARDISPMODE[2], _6I4446_$1I3863_TXCHARDISPMODE_2__vlIN);
 reg [1:16] _6I4446_$1I3863_TXCHARDISPMODE_1__vlIN;
 cstw cstw_587_1 (_6I4446_$1I3863_TXCHARDISPMODE[1], _6I4446_$1I3863_TXCHARDISPMODE_1__vlIN);
 reg [1:16] _6I4446_$1I3863_TXCHARDISPMODE_0__vlIN;
 cstw cstw_587_0 (_6I4446_$1I3863_TXCHARDISPMODE[0], _6I4446_$1I3863_TXCHARDISPMODE_0__vlIN);

 wire [3:0] _6I4446_$1I3863_TXCHARDISPVAL;
 reg [1:16] _6I4446_$1I3863_TXCHARDISPVAL_3__vlIN;
 cstw cstw_588_3 (_6I4446_$1I3863_TXCHARDISPVAL[3], _6I4446_$1I3863_TXCHARDISPVAL_3__vlIN);
 reg [1:16] _6I4446_$1I3863_TXCHARDISPVAL_2__vlIN;
 cstw cstw_588_2 (_6I4446_$1I3863_TXCHARDISPVAL[2], _6I4446_$1I3863_TXCHARDISPVAL_2__vlIN);
 reg [1:16] _6I4446_$1I3863_TXCHARDISPVAL_1__vlIN;
 cstw cstw_588_1 (_6I4446_$1I3863_TXCHARDISPVAL[1], _6I4446_$1I3863_TXCHARDISPVAL_1__vlIN);
 reg [1:16] _6I4446_$1I3863_TXCHARDISPVAL_0__vlIN;
 cstw cstw_588_0 (_6I4446_$1I3863_TXCHARDISPVAL[0], _6I4446_$1I3863_TXCHARDISPVAL_0__vlIN);

 wire [3:0] _6I4446_$1I3863_TXCHARISK;
 reg [1:16] _6I4446_$1I3863_TXCHARISK_3__vlIN;
 cstw cstw_589_3 (_6I4446_$1I3863_TXCHARISK[3], _6I4446_$1I3863_TXCHARISK_3__vlIN);
 reg [1:16] _6I4446_$1I3863_TXCHARISK_2__vlIN;
 cstw cstw_589_2 (_6I4446_$1I3863_TXCHARISK[2], _6I4446_$1I3863_TXCHARISK_2__vlIN);
 reg [1:16] _6I4446_$1I3863_TXCHARISK_1__vlIN;
 cstw cstw_589_1 (_6I4446_$1I3863_TXCHARISK[1], _6I4446_$1I3863_TXCHARISK_1__vlIN);
 reg [1:16] _6I4446_$1I3863_TXCHARISK_0__vlIN;
 cstw cstw_589_0 (_6I4446_$1I3863_TXCHARISK[0], _6I4446_$1I3863_TXCHARISK_0__vlIN);

 wire [31:0] _6I4446_$1I3863_TXDATA;
 reg [1:16] _6I4446_$1I3863_TXDATA_31__vlIN;
 cstw cstw_590_31 (_6I4446_$1I3863_TXDATA[31], _6I4446_$1I3863_TXDATA_31__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_30__vlIN;
 cstw cstw_590_30 (_6I4446_$1I3863_TXDATA[30], _6I4446_$1I3863_TXDATA_30__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_29__vlIN;
 cstw cstw_590_29 (_6I4446_$1I3863_TXDATA[29], _6I4446_$1I3863_TXDATA_29__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_28__vlIN;
 cstw cstw_590_28 (_6I4446_$1I3863_TXDATA[28], _6I4446_$1I3863_TXDATA_28__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_27__vlIN;
 cstw cstw_590_27 (_6I4446_$1I3863_TXDATA[27], _6I4446_$1I3863_TXDATA_27__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_26__vlIN;
 cstw cstw_590_26 (_6I4446_$1I3863_TXDATA[26], _6I4446_$1I3863_TXDATA_26__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_25__vlIN;
 cstw cstw_590_25 (_6I4446_$1I3863_TXDATA[25], _6I4446_$1I3863_TXDATA_25__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_24__vlIN;
 cstw cstw_590_24 (_6I4446_$1I3863_TXDATA[24], _6I4446_$1I3863_TXDATA_24__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_23__vlIN;
 cstw cstw_590_23 (_6I4446_$1I3863_TXDATA[23], _6I4446_$1I3863_TXDATA_23__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_22__vlIN;
 cstw cstw_590_22 (_6I4446_$1I3863_TXDATA[22], _6I4446_$1I3863_TXDATA_22__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_21__vlIN;
 cstw cstw_590_21 (_6I4446_$1I3863_TXDATA[21], _6I4446_$1I3863_TXDATA_21__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_20__vlIN;
 cstw cstw_590_20 (_6I4446_$1I3863_TXDATA[20], _6I4446_$1I3863_TXDATA_20__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_19__vlIN;
 cstw cstw_590_19 (_6I4446_$1I3863_TXDATA[19], _6I4446_$1I3863_TXDATA_19__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_18__vlIN;
 cstw cstw_590_18 (_6I4446_$1I3863_TXDATA[18], _6I4446_$1I3863_TXDATA_18__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_17__vlIN;
 cstw cstw_590_17 (_6I4446_$1I3863_TXDATA[17], _6I4446_$1I3863_TXDATA_17__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_16__vlIN;
 cstw cstw_590_16 (_6I4446_$1I3863_TXDATA[16], _6I4446_$1I3863_TXDATA_16__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_15__vlIN;
 cstw cstw_590_15 (_6I4446_$1I3863_TXDATA[15], _6I4446_$1I3863_TXDATA_15__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_14__vlIN;
 cstw cstw_590_14 (_6I4446_$1I3863_TXDATA[14], _6I4446_$1I3863_TXDATA_14__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_13__vlIN;
 cstw cstw_590_13 (_6I4446_$1I3863_TXDATA[13], _6I4446_$1I3863_TXDATA_13__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_12__vlIN;
 cstw cstw_590_12 (_6I4446_$1I3863_TXDATA[12], _6I4446_$1I3863_TXDATA_12__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_11__vlIN;
 cstw cstw_590_11 (_6I4446_$1I3863_TXDATA[11], _6I4446_$1I3863_TXDATA_11__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_10__vlIN;
 cstw cstw_590_10 (_6I4446_$1I3863_TXDATA[10], _6I4446_$1I3863_TXDATA_10__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_9__vlIN;
 cstw cstw_590_9 (_6I4446_$1I3863_TXDATA[9], _6I4446_$1I3863_TXDATA_9__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_8__vlIN;
 cstw cstw_590_8 (_6I4446_$1I3863_TXDATA[8], _6I4446_$1I3863_TXDATA_8__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_7__vlIN;
 cstw cstw_590_7 (_6I4446_$1I3863_TXDATA[7], _6I4446_$1I3863_TXDATA_7__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_6__vlIN;
 cstw cstw_590_6 (_6I4446_$1I3863_TXDATA[6], _6I4446_$1I3863_TXDATA_6__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_5__vlIN;
 cstw cstw_590_5 (_6I4446_$1I3863_TXDATA[5], _6I4446_$1I3863_TXDATA_5__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_4__vlIN;
 cstw cstw_590_4 (_6I4446_$1I3863_TXDATA[4], _6I4446_$1I3863_TXDATA_4__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_3__vlIN;
 cstw cstw_590_3 (_6I4446_$1I3863_TXDATA[3], _6I4446_$1I3863_TXDATA_3__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_2__vlIN;
 cstw cstw_590_2 (_6I4446_$1I3863_TXDATA[2], _6I4446_$1I3863_TXDATA_2__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_1__vlIN;
 cstw cstw_590_1 (_6I4446_$1I3863_TXDATA[1], _6I4446_$1I3863_TXDATA_1__vlIN);
 reg [1:16] _6I4446_$1I3863_TXDATA_0__vlIN;
 cstw cstw_590_0 (_6I4446_$1I3863_TXDATA[0], _6I4446_$1I3863_TXDATA_0__vlIN);

 wire  _6I4446_$1I3863_TXFORCECRCERR;
 reg [1:16] _6I4446_$1I3863_TXFORCECRCERR__vlIN;
 cstw cstw_591 (_6I4446_$1I3863_TXFORCECRCERR, _6I4446_$1I3863_TXFORCECRCERR__vlIN);

 wire  _6I4446_$1I3863_TXINHIBIT;
 reg [1:16] _6I4446_$1I3863_TXINHIBIT__vlIN;
 cstw cstw_592 (_6I4446_$1I3863_TXINHIBIT, _6I4446_$1I3863_TXINHIBIT__vlIN);

 wire  _6I4446_$1I3863_TXPOLARITY;
 reg [1:16] _6I4446_$1I3863_TXPOLARITY__vlIN;
 cstw cstw_593 (_6I4446_$1I3863_TXPOLARITY, _6I4446_$1I3863_TXPOLARITY__vlIN);

 wire  _6I4446_$1I3863_TXRESET;
 reg [1:16] _6I4446_$1I3863_TXRESET__vlIN;
 cstw cstw_594 (_6I4446_$1I3863_TXRESET, _6I4446_$1I3863_TXRESET__vlIN);

 wire  _6I4446_$1I3863_TXUSRCLK;
 reg [1:16] _6I4446_$1I3863_TXUSRCLK__vlIN;
 cstw cstw_595 (_6I4446_$1I3863_TXUSRCLK, _6I4446_$1I3863_TXUSRCLK__vlIN);

 wire  _6I4446_$1I3863_TXUSRCLK2;
 reg [1:16] _6I4446_$1I3863_TXUSRCLK2__vlIN;
 cstw cstw_596 (_6I4446_$1I3863_TXUSRCLK2, _6I4446_$1I3863_TXUSRCLK2__vlIN);

 GT_CUSTOM _6I4446_$1I3863 ( _6I4446_$1I3863_CHBONDDONE , _6I4446_$1I3863_CHBONDO , _6I4446_$1I3863_CONFIGOUT , _6I4446_$1I3863_RXBUFSTATUS , _6I4446_$1I3863_RXCHARISCOMMA , _6I4446_$1I3863_RXCHARISK , _6I4446_$1I3863_RXCHECKINGCRC , _6I4446_$1I3863_RXCLKCORCNT , _6I4446_$1I3863_RXCOMMADET , _6I4446_$1I3863_RXCRCERR , _6I4446_$1I3863_RXDATA , _6I4446_$1I3863_RXDISPERR , _6I4446_$1I3863_RXLOSSOFSYNC , _6I4446_$1I3863_RXNOTINTABLE , _6I4446_$1I3863_RXREALIGN , _6I4446_$1I3863_RXRECCLK , _6I4446_$1I3863_RXRUNDISP , _6I4446_$1I3863_TXBUFERR , _6I4446_$1I3863_TXKERR , _6I4446_$1I3863_TXN , _6I4446_$1I3863_TXP , _6I4446_$1I3863_TXRUNDISP , _6I4446_$1I3863_BREFCLK , _6I4446_$1I3863_BREFCLK2 , _6I4446_$1I3863_CHBONDI , _6I4446_$1I3863_CONFIGENABLE , _6I4446_$1I3863_CONFIGIN , _6I4446_$1I3863_ENCHANSYNC , _6I4446_$1I3863_ENMCOMMAALIGN , _6I4446_$1I3863_ENPCOMMAALIGN , _6I4446_$1I3863_LOOPBACK , _6I4446_$1I3863_POWERDOWN , _6I4446_$1I3863_REFCLK , _6I4446_$1I3863_REFCLK2 , _6I4446_$1I3863_REFCLKSEL , _6I4446_$1I3863_RXN , _6I4446_$1I3863_RXP , _6I4446_$1I3863_RXPOLARITY , _6I4446_$1I3863_RXRESET , _6I4446_$1I3863_RXUSRCLK , _6I4446_$1I3863_RXUSRCLK2 , _6I4446_$1I3863_TXBYPASS8B10B , _6I4446_$1I3863_TXCHARDISPMODE , _6I4446_$1I3863_TXCHARDISPVAL , _6I4446_$1I3863_TXCHARISK , _6I4446_$1I3863_TXDATA , _6I4446_$1I3863_TXFORCECRCERR , _6I4446_$1I3863_TXINHIBIT , _6I4446_$1I3863_TXPOLARITY , _6I4446_$1I3863_TXRESET , _6I4446_$1I3863_TXUSRCLK , _6I4446_$1I3863_TXUSRCLK2  );

// ----------------------------------- //

 wire [4:0] _6I4415_$1I4152_din;
 reg [1:16] _6I4415_$1I4152_din_4__vlIN;
 cstw cstw_597_4 (_6I4415_$1I4152_din[4], _6I4415_$1I4152_din_4__vlIN);
 reg [1:16] _6I4415_$1I4152_din_3__vlIN;
 cstw cstw_597_3 (_6I4415_$1I4152_din[3], _6I4415_$1I4152_din_3__vlIN);
 reg [1:16] _6I4415_$1I4152_din_2__vlIN;
 cstw cstw_597_2 (_6I4415_$1I4152_din[2], _6I4415_$1I4152_din_2__vlIN);
 reg [1:16] _6I4415_$1I4152_din_1__vlIN;
 cstw cstw_597_1 (_6I4415_$1I4152_din[1], _6I4415_$1I4152_din_1__vlIN);
 reg [1:16] _6I4415_$1I4152_din_0__vlIN;
 cstw cstw_597_0 (_6I4415_$1I4152_din[0], _6I4415_$1I4152_din_0__vlIN);

 wire  _6I4415_$1I4152_wr_en;
 reg [1:16] _6I4415_$1I4152_wr_en__vlIN;
 cstw cstw_598 (_6I4415_$1I4152_wr_en, _6I4415_$1I4152_wr_en__vlIN);

 wire  _6I4415_$1I4152_wr_clk;
 reg [1:16] _6I4415_$1I4152_wr_clk__vlIN;
 cstw cstw_599 (_6I4415_$1I4152_wr_clk, _6I4415_$1I4152_wr_clk__vlIN);

 wire  _6I4415_$1I4152_rd_en;
 reg [1:16] _6I4415_$1I4152_rd_en__vlIN;
 cstw cstw_600 (_6I4415_$1I4152_rd_en, _6I4415_$1I4152_rd_en__vlIN);

 wire  _6I4415_$1I4152_rd_clk;
 reg [1:16] _6I4415_$1I4152_rd_clk__vlIN;
 cstw cstw_601 (_6I4415_$1I4152_rd_clk, _6I4415_$1I4152_rd_clk__vlIN);

 wire  _6I4415_$1I4152_ainit;
 reg [1:16] _6I4415_$1I4152_ainit__vlIN;
 cstw cstw_602 (_6I4415_$1I4152_ainit, _6I4415_$1I4152_ainit__vlIN);

 wire [4:0] _6I4415_$1I4152_dout;

 wire  _6I4415_$1I4152_full;

 wire  _6I4415_$1I4152_empty;

 af_clb_5x31rpm _6I4415_$1I4152 ( _6I4415_$1I4152_din , _6I4415_$1I4152_wr_en , _6I4415_$1I4152_wr_clk , _6I4415_$1I4152_rd_en , _6I4415_$1I4152_rd_clk , _6I4415_$1I4152_ainit , _6I4415_$1I4152_dout , _6I4415_$1I4152_full , _6I4415_$1I4152_empty  );

// ----------------------------------- //

 wire  _6I4415_$1I3863_CHBONDDONE;

 wire [3:0] _6I4415_$1I3863_CHBONDO;

 wire  _6I4415_$1I3863_CONFIGOUT;

 wire [1:0] _6I4415_$1I3863_RXBUFSTATUS;

 wire [3:0] _6I4415_$1I3863_RXCHARISCOMMA;

 wire [3:0] _6I4415_$1I3863_RXCHARISK;

 wire  _6I4415_$1I3863_RXCHECKINGCRC;

 wire [2:0] _6I4415_$1I3863_RXCLKCORCNT;

 wire  _6I4415_$1I3863_RXCOMMADET;

 wire  _6I4415_$1I3863_RXCRCERR;

 wire [31:0] _6I4415_$1I3863_RXDATA;

 wire [3:0] _6I4415_$1I3863_RXDISPERR;

 wire [1:0] _6I4415_$1I3863_RXLOSSOFSYNC;

 wire [3:0] _6I4415_$1I3863_RXNOTINTABLE;

 wire  _6I4415_$1I3863_RXREALIGN;

 wire  _6I4415_$1I3863_RXRECCLK;

 wire [3:0] _6I4415_$1I3863_RXRUNDISP;

 wire  _6I4415_$1I3863_TXBUFERR;

 wire [3:0] _6I4415_$1I3863_TXKERR;

 wire  _6I4415_$1I3863_TXN;

 wire  _6I4415_$1I3863_TXP;

 wire [3:0] _6I4415_$1I3863_TXRUNDISP;

 wire  _6I4415_$1I3863_BREFCLK;
 reg [1:16] _6I4415_$1I3863_BREFCLK__vlIN;
 cstw cstw_603 (_6I4415_$1I3863_BREFCLK, _6I4415_$1I3863_BREFCLK__vlIN);

 wire  _6I4415_$1I3863_BREFCLK2;
 reg [1:16] _6I4415_$1I3863_BREFCLK2__vlIN;
 cstw cstw_604 (_6I4415_$1I3863_BREFCLK2, _6I4415_$1I3863_BREFCLK2__vlIN);

 wire [3:0] _6I4415_$1I3863_CHBONDI;
 reg [1:16] _6I4415_$1I3863_CHBONDI_3__vlIN;
 cstw cstw_605_3 (_6I4415_$1I3863_CHBONDI[3], _6I4415_$1I3863_CHBONDI_3__vlIN);
 reg [1:16] _6I4415_$1I3863_CHBONDI_2__vlIN;
 cstw cstw_605_2 (_6I4415_$1I3863_CHBONDI[2], _6I4415_$1I3863_CHBONDI_2__vlIN);
 reg [1:16] _6I4415_$1I3863_CHBONDI_1__vlIN;
 cstw cstw_605_1 (_6I4415_$1I3863_CHBONDI[1], _6I4415_$1I3863_CHBONDI_1__vlIN);
 reg [1:16] _6I4415_$1I3863_CHBONDI_0__vlIN;
 cstw cstw_605_0 (_6I4415_$1I3863_CHBONDI[0], _6I4415_$1I3863_CHBONDI_0__vlIN);

 wire  _6I4415_$1I3863_CONFIGENABLE;
 reg [1:16] _6I4415_$1I3863_CONFIGENABLE__vlIN;
 cstw cstw_606 (_6I4415_$1I3863_CONFIGENABLE, _6I4415_$1I3863_CONFIGENABLE__vlIN);

 wire  _6I4415_$1I3863_CONFIGIN;
 reg [1:16] _6I4415_$1I3863_CONFIGIN__vlIN;
 cstw cstw_607 (_6I4415_$1I3863_CONFIGIN, _6I4415_$1I3863_CONFIGIN__vlIN);

 wire  _6I4415_$1I3863_ENCHANSYNC;
 reg [1:16] _6I4415_$1I3863_ENCHANSYNC__vlIN;
 cstw cstw_608 (_6I4415_$1I3863_ENCHANSYNC, _6I4415_$1I3863_ENCHANSYNC__vlIN);

 wire  _6I4415_$1I3863_ENMCOMMAALIGN;
 reg [1:16] _6I4415_$1I3863_ENMCOMMAALIGN__vlIN;
 cstw cstw_609 (_6I4415_$1I3863_ENMCOMMAALIGN, _6I4415_$1I3863_ENMCOMMAALIGN__vlIN);

 wire  _6I4415_$1I3863_ENPCOMMAALIGN;
 reg [1:16] _6I4415_$1I3863_ENPCOMMAALIGN__vlIN;
 cstw cstw_610 (_6I4415_$1I3863_ENPCOMMAALIGN, _6I4415_$1I3863_ENPCOMMAALIGN__vlIN);

 wire [1:0] _6I4415_$1I3863_LOOPBACK;
 reg [1:16] _6I4415_$1I3863_LOOPBACK_1__vlIN;
 cstw cstw_611_1 (_6I4415_$1I3863_LOOPBACK[1], _6I4415_$1I3863_LOOPBACK_1__vlIN);
 reg [1:16] _6I4415_$1I3863_LOOPBACK_0__vlIN;
 cstw cstw_611_0 (_6I4415_$1I3863_LOOPBACK[0], _6I4415_$1I3863_LOOPBACK_0__vlIN);

 wire  _6I4415_$1I3863_POWERDOWN;
 reg [1:16] _6I4415_$1I3863_POWERDOWN__vlIN;
 cstw cstw_612 (_6I4415_$1I3863_POWERDOWN, _6I4415_$1I3863_POWERDOWN__vlIN);

 wire  _6I4415_$1I3863_REFCLK;
 reg [1:16] _6I4415_$1I3863_REFCLK__vlIN;
 cstw cstw_613 (_6I4415_$1I3863_REFCLK, _6I4415_$1I3863_REFCLK__vlIN);

 wire  _6I4415_$1I3863_REFCLK2;
 reg [1:16] _6I4415_$1I3863_REFCLK2__vlIN;
 cstw cstw_614 (_6I4415_$1I3863_REFCLK2, _6I4415_$1I3863_REFCLK2__vlIN);

 wire  _6I4415_$1I3863_REFCLKSEL;
 reg [1:16] _6I4415_$1I3863_REFCLKSEL__vlIN;
 cstw cstw_615 (_6I4415_$1I3863_REFCLKSEL, _6I4415_$1I3863_REFCLKSEL__vlIN);

 wire  _6I4415_$1I3863_RXN;
 reg [1:16] _6I4415_$1I3863_RXN__vlIN;
 cstw cstw_616 (_6I4415_$1I3863_RXN, _6I4415_$1I3863_RXN__vlIN);

 wire  _6I4415_$1I3863_RXP;
 reg [1:16] _6I4415_$1I3863_RXP__vlIN;
 cstw cstw_617 (_6I4415_$1I3863_RXP, _6I4415_$1I3863_RXP__vlIN);

 wire  _6I4415_$1I3863_RXPOLARITY;
 reg [1:16] _6I4415_$1I3863_RXPOLARITY__vlIN;
 cstw cstw_618 (_6I4415_$1I3863_RXPOLARITY, _6I4415_$1I3863_RXPOLARITY__vlIN);

 wire  _6I4415_$1I3863_RXRESET;
 reg [1:16] _6I4415_$1I3863_RXRESET__vlIN;
 cstw cstw_619 (_6I4415_$1I3863_RXRESET, _6I4415_$1I3863_RXRESET__vlIN);

 wire  _6I4415_$1I3863_RXUSRCLK;
 reg [1:16] _6I4415_$1I3863_RXUSRCLK__vlIN;
 cstw cstw_620 (_6I4415_$1I3863_RXUSRCLK, _6I4415_$1I3863_RXUSRCLK__vlIN);

 wire  _6I4415_$1I3863_RXUSRCLK2;
 reg [1:16] _6I4415_$1I3863_RXUSRCLK2__vlIN;
 cstw cstw_621 (_6I4415_$1I3863_RXUSRCLK2, _6I4415_$1I3863_RXUSRCLK2__vlIN);

 wire [3:0] _6I4415_$1I3863_TXBYPASS8B10B;
 reg [1:16] _6I4415_$1I3863_TXBYPASS8B10B_3__vlIN;
 cstw cstw_622_3 (_6I4415_$1I3863_TXBYPASS8B10B[3], _6I4415_$1I3863_TXBYPASS8B10B_3__vlIN);
 reg [1:16] _6I4415_$1I3863_TXBYPASS8B10B_2__vlIN;
 cstw cstw_622_2 (_6I4415_$1I3863_TXBYPASS8B10B[2], _6I4415_$1I3863_TXBYPASS8B10B_2__vlIN);
 reg [1:16] _6I4415_$1I3863_TXBYPASS8B10B_1__vlIN;
 cstw cstw_622_1 (_6I4415_$1I3863_TXBYPASS8B10B[1], _6I4415_$1I3863_TXBYPASS8B10B_1__vlIN);
 reg [1:16] _6I4415_$1I3863_TXBYPASS8B10B_0__vlIN;
 cstw cstw_622_0 (_6I4415_$1I3863_TXBYPASS8B10B[0], _6I4415_$1I3863_TXBYPASS8B10B_0__vlIN);

 wire [3:0] _6I4415_$1I3863_TXCHARDISPMODE;
 reg [1:16] _6I4415_$1I3863_TXCHARDISPMODE_3__vlIN;
 cstw cstw_623_3 (_6I4415_$1I3863_TXCHARDISPMODE[3], _6I4415_$1I3863_TXCHARDISPMODE_3__vlIN);
 reg [1:16] _6I4415_$1I3863_TXCHARDISPMODE_2__vlIN;
 cstw cstw_623_2 (_6I4415_$1I3863_TXCHARDISPMODE[2], _6I4415_$1I3863_TXCHARDISPMODE_2__vlIN);
 reg [1:16] _6I4415_$1I3863_TXCHARDISPMODE_1__vlIN;
 cstw cstw_623_1 (_6I4415_$1I3863_TXCHARDISPMODE[1], _6I4415_$1I3863_TXCHARDISPMODE_1__vlIN);
 reg [1:16] _6I4415_$1I3863_TXCHARDISPMODE_0__vlIN;
 cstw cstw_623_0 (_6I4415_$1I3863_TXCHARDISPMODE[0], _6I4415_$1I3863_TXCHARDISPMODE_0__vlIN);

 wire [3:0] _6I4415_$1I3863_TXCHARDISPVAL;
 reg [1:16] _6I4415_$1I3863_TXCHARDISPVAL_3__vlIN;
 cstw cstw_624_3 (_6I4415_$1I3863_TXCHARDISPVAL[3], _6I4415_$1I3863_TXCHARDISPVAL_3__vlIN);
 reg [1:16] _6I4415_$1I3863_TXCHARDISPVAL_2__vlIN;
 cstw cstw_624_2 (_6I4415_$1I3863_TXCHARDISPVAL[2], _6I4415_$1I3863_TXCHARDISPVAL_2__vlIN);
 reg [1:16] _6I4415_$1I3863_TXCHARDISPVAL_1__vlIN;
 cstw cstw_624_1 (_6I4415_$1I3863_TXCHARDISPVAL[1], _6I4415_$1I3863_TXCHARDISPVAL_1__vlIN);
 reg [1:16] _6I4415_$1I3863_TXCHARDISPVAL_0__vlIN;
 cstw cstw_624_0 (_6I4415_$1I3863_TXCHARDISPVAL[0], _6I4415_$1I3863_TXCHARDISPVAL_0__vlIN);

 wire [3:0] _6I4415_$1I3863_TXCHARISK;
 reg [1:16] _6I4415_$1I3863_TXCHARISK_3__vlIN;
 cstw cstw_625_3 (_6I4415_$1I3863_TXCHARISK[3], _6I4415_$1I3863_TXCHARISK_3__vlIN);
 reg [1:16] _6I4415_$1I3863_TXCHARISK_2__vlIN;
 cstw cstw_625_2 (_6I4415_$1I3863_TXCHARISK[2], _6I4415_$1I3863_TXCHARISK_2__vlIN);
 reg [1:16] _6I4415_$1I3863_TXCHARISK_1__vlIN;
 cstw cstw_625_1 (_6I4415_$1I3863_TXCHARISK[1], _6I4415_$1I3863_TXCHARISK_1__vlIN);
 reg [1:16] _6I4415_$1I3863_TXCHARISK_0__vlIN;
 cstw cstw_625_0 (_6I4415_$1I3863_TXCHARISK[0], _6I4415_$1I3863_TXCHARISK_0__vlIN);

 wire [31:0] _6I4415_$1I3863_TXDATA;
 reg [1:16] _6I4415_$1I3863_TXDATA_31__vlIN;
 cstw cstw_626_31 (_6I4415_$1I3863_TXDATA[31], _6I4415_$1I3863_TXDATA_31__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_30__vlIN;
 cstw cstw_626_30 (_6I4415_$1I3863_TXDATA[30], _6I4415_$1I3863_TXDATA_30__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_29__vlIN;
 cstw cstw_626_29 (_6I4415_$1I3863_TXDATA[29], _6I4415_$1I3863_TXDATA_29__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_28__vlIN;
 cstw cstw_626_28 (_6I4415_$1I3863_TXDATA[28], _6I4415_$1I3863_TXDATA_28__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_27__vlIN;
 cstw cstw_626_27 (_6I4415_$1I3863_TXDATA[27], _6I4415_$1I3863_TXDATA_27__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_26__vlIN;
 cstw cstw_626_26 (_6I4415_$1I3863_TXDATA[26], _6I4415_$1I3863_TXDATA_26__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_25__vlIN;
 cstw cstw_626_25 (_6I4415_$1I3863_TXDATA[25], _6I4415_$1I3863_TXDATA_25__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_24__vlIN;
 cstw cstw_626_24 (_6I4415_$1I3863_TXDATA[24], _6I4415_$1I3863_TXDATA_24__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_23__vlIN;
 cstw cstw_626_23 (_6I4415_$1I3863_TXDATA[23], _6I4415_$1I3863_TXDATA_23__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_22__vlIN;
 cstw cstw_626_22 (_6I4415_$1I3863_TXDATA[22], _6I4415_$1I3863_TXDATA_22__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_21__vlIN;
 cstw cstw_626_21 (_6I4415_$1I3863_TXDATA[21], _6I4415_$1I3863_TXDATA_21__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_20__vlIN;
 cstw cstw_626_20 (_6I4415_$1I3863_TXDATA[20], _6I4415_$1I3863_TXDATA_20__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_19__vlIN;
 cstw cstw_626_19 (_6I4415_$1I3863_TXDATA[19], _6I4415_$1I3863_TXDATA_19__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_18__vlIN;
 cstw cstw_626_18 (_6I4415_$1I3863_TXDATA[18], _6I4415_$1I3863_TXDATA_18__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_17__vlIN;
 cstw cstw_626_17 (_6I4415_$1I3863_TXDATA[17], _6I4415_$1I3863_TXDATA_17__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_16__vlIN;
 cstw cstw_626_16 (_6I4415_$1I3863_TXDATA[16], _6I4415_$1I3863_TXDATA_16__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_15__vlIN;
 cstw cstw_626_15 (_6I4415_$1I3863_TXDATA[15], _6I4415_$1I3863_TXDATA_15__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_14__vlIN;
 cstw cstw_626_14 (_6I4415_$1I3863_TXDATA[14], _6I4415_$1I3863_TXDATA_14__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_13__vlIN;
 cstw cstw_626_13 (_6I4415_$1I3863_TXDATA[13], _6I4415_$1I3863_TXDATA_13__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_12__vlIN;
 cstw cstw_626_12 (_6I4415_$1I3863_TXDATA[12], _6I4415_$1I3863_TXDATA_12__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_11__vlIN;
 cstw cstw_626_11 (_6I4415_$1I3863_TXDATA[11], _6I4415_$1I3863_TXDATA_11__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_10__vlIN;
 cstw cstw_626_10 (_6I4415_$1I3863_TXDATA[10], _6I4415_$1I3863_TXDATA_10__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_9__vlIN;
 cstw cstw_626_9 (_6I4415_$1I3863_TXDATA[9], _6I4415_$1I3863_TXDATA_9__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_8__vlIN;
 cstw cstw_626_8 (_6I4415_$1I3863_TXDATA[8], _6I4415_$1I3863_TXDATA_8__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_7__vlIN;
 cstw cstw_626_7 (_6I4415_$1I3863_TXDATA[7], _6I4415_$1I3863_TXDATA_7__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_6__vlIN;
 cstw cstw_626_6 (_6I4415_$1I3863_TXDATA[6], _6I4415_$1I3863_TXDATA_6__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_5__vlIN;
 cstw cstw_626_5 (_6I4415_$1I3863_TXDATA[5], _6I4415_$1I3863_TXDATA_5__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_4__vlIN;
 cstw cstw_626_4 (_6I4415_$1I3863_TXDATA[4], _6I4415_$1I3863_TXDATA_4__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_3__vlIN;
 cstw cstw_626_3 (_6I4415_$1I3863_TXDATA[3], _6I4415_$1I3863_TXDATA_3__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_2__vlIN;
 cstw cstw_626_2 (_6I4415_$1I3863_TXDATA[2], _6I4415_$1I3863_TXDATA_2__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_1__vlIN;
 cstw cstw_626_1 (_6I4415_$1I3863_TXDATA[1], _6I4415_$1I3863_TXDATA_1__vlIN);
 reg [1:16] _6I4415_$1I3863_TXDATA_0__vlIN;
 cstw cstw_626_0 (_6I4415_$1I3863_TXDATA[0], _6I4415_$1I3863_TXDATA_0__vlIN);

 wire  _6I4415_$1I3863_TXFORCECRCERR;
 reg [1:16] _6I4415_$1I3863_TXFORCECRCERR__vlIN;
 cstw cstw_627 (_6I4415_$1I3863_TXFORCECRCERR, _6I4415_$1I3863_TXFORCECRCERR__vlIN);

 wire  _6I4415_$1I3863_TXINHIBIT;
 reg [1:16] _6I4415_$1I3863_TXINHIBIT__vlIN;
 cstw cstw_628 (_6I4415_$1I3863_TXINHIBIT, _6I4415_$1I3863_TXINHIBIT__vlIN);

 wire  _6I4415_$1I3863_TXPOLARITY;
 reg [1:16] _6I4415_$1I3863_TXPOLARITY__vlIN;
 cstw cstw_629 (_6I4415_$1I3863_TXPOLARITY, _6I4415_$1I3863_TXPOLARITY__vlIN);

 wire  _6I4415_$1I3863_TXRESET;
 reg [1:16] _6I4415_$1I3863_TXRESET__vlIN;
 cstw cstw_630 (_6I4415_$1I3863_TXRESET, _6I4415_$1I3863_TXRESET__vlIN);

 wire  _6I4415_$1I3863_TXUSRCLK;
 reg [1:16] _6I4415_$1I3863_TXUSRCLK__vlIN;
 cstw cstw_631 (_6I4415_$1I3863_TXUSRCLK, _6I4415_$1I3863_TXUSRCLK__vlIN);

 wire  _6I4415_$1I3863_TXUSRCLK2;
 reg [1:16] _6I4415_$1I3863_TXUSRCLK2__vlIN;
 cstw cstw_632 (_6I4415_$1I3863_TXUSRCLK2, _6I4415_$1I3863_TXUSRCLK2__vlIN);

 GT_CUSTOM _6I4415_$1I3863 ( _6I4415_$1I3863_CHBONDDONE , _6I4415_$1I3863_CHBONDO , _6I4415_$1I3863_CONFIGOUT , _6I4415_$1I3863_RXBUFSTATUS , _6I4415_$1I3863_RXCHARISCOMMA , _6I4415_$1I3863_RXCHARISK , _6I4415_$1I3863_RXCHECKINGCRC , _6I4415_$1I3863_RXCLKCORCNT , _6I4415_$1I3863_RXCOMMADET , _6I4415_$1I3863_RXCRCERR , _6I4415_$1I3863_RXDATA , _6I4415_$1I3863_RXDISPERR , _6I4415_$1I3863_RXLOSSOFSYNC , _6I4415_$1I3863_RXNOTINTABLE , _6I4415_$1I3863_RXREALIGN , _6I4415_$1I3863_RXRECCLK , _6I4415_$1I3863_RXRUNDISP , _6I4415_$1I3863_TXBUFERR , _6I4415_$1I3863_TXKERR , _6I4415_$1I3863_TXN , _6I4415_$1I3863_TXP , _6I4415_$1I3863_TXRUNDISP , _6I4415_$1I3863_BREFCLK , _6I4415_$1I3863_BREFCLK2 , _6I4415_$1I3863_CHBONDI , _6I4415_$1I3863_CONFIGENABLE , _6I4415_$1I3863_CONFIGIN , _6I4415_$1I3863_ENCHANSYNC , _6I4415_$1I3863_ENMCOMMAALIGN , _6I4415_$1I3863_ENPCOMMAALIGN , _6I4415_$1I3863_LOOPBACK , _6I4415_$1I3863_POWERDOWN , _6I4415_$1I3863_REFCLK , _6I4415_$1I3863_REFCLK2 , _6I4415_$1I3863_REFCLKSEL , _6I4415_$1I3863_RXN , _6I4415_$1I3863_RXP , _6I4415_$1I3863_RXPOLARITY , _6I4415_$1I3863_RXRESET , _6I4415_$1I3863_RXUSRCLK , _6I4415_$1I3863_RXUSRCLK2 , _6I4415_$1I3863_TXBYPASS8B10B , _6I4415_$1I3863_TXCHARDISPMODE , _6I4415_$1I3863_TXCHARDISPVAL , _6I4415_$1I3863_TXCHARISK , _6I4415_$1I3863_TXDATA , _6I4415_$1I3863_TXFORCECRCERR , _6I4415_$1I3863_TXINHIBIT , _6I4415_$1I3863_TXPOLARITY , _6I4415_$1I3863_TXRESET , _6I4415_$1I3863_TXUSRCLK , _6I4415_$1I3863_TXUSRCLK2  );

// ----------------------------------- //

 wire [4:0] _6I4412_$1I4152_din;
 reg [1:16] _6I4412_$1I4152_din_4__vlIN;
 cstw cstw_633_4 (_6I4412_$1I4152_din[4], _6I4412_$1I4152_din_4__vlIN);
 reg [1:16] _6I4412_$1I4152_din_3__vlIN;
 cstw cstw_633_3 (_6I4412_$1I4152_din[3], _6I4412_$1I4152_din_3__vlIN);
 reg [1:16] _6I4412_$1I4152_din_2__vlIN;
 cstw cstw_633_2 (_6I4412_$1I4152_din[2], _6I4412_$1I4152_din_2__vlIN);
 reg [1:16] _6I4412_$1I4152_din_1__vlIN;
 cstw cstw_633_1 (_6I4412_$1I4152_din[1], _6I4412_$1I4152_din_1__vlIN);
 reg [1:16] _6I4412_$1I4152_din_0__vlIN;
 cstw cstw_633_0 (_6I4412_$1I4152_din[0], _6I4412_$1I4152_din_0__vlIN);

 wire  _6I4412_$1I4152_wr_en;
 reg [1:16] _6I4412_$1I4152_wr_en__vlIN;
 cstw cstw_634 (_6I4412_$1I4152_wr_en, _6I4412_$1I4152_wr_en__vlIN);

 wire  _6I4412_$1I4152_wr_clk;
 reg [1:16] _6I4412_$1I4152_wr_clk__vlIN;
 cstw cstw_635 (_6I4412_$1I4152_wr_clk, _6I4412_$1I4152_wr_clk__vlIN);

 wire  _6I4412_$1I4152_rd_en;
 reg [1:16] _6I4412_$1I4152_rd_en__vlIN;
 cstw cstw_636 (_6I4412_$1I4152_rd_en, _6I4412_$1I4152_rd_en__vlIN);

 wire  _6I4412_$1I4152_rd_clk;
 reg [1:16] _6I4412_$1I4152_rd_clk__vlIN;
 cstw cstw_637 (_6I4412_$1I4152_rd_clk, _6I4412_$1I4152_rd_clk__vlIN);

 wire  _6I4412_$1I4152_ainit;
 reg [1:16] _6I4412_$1I4152_ainit__vlIN;
 cstw cstw_638 (_6I4412_$1I4152_ainit, _6I4412_$1I4152_ainit__vlIN);

 wire [4:0] _6I4412_$1I4152_dout;

 wire  _6I4412_$1I4152_full;

 wire  _6I4412_$1I4152_empty;

 af_clb_5x31rpm _6I4412_$1I4152 ( _6I4412_$1I4152_din , _6I4412_$1I4152_wr_en , _6I4412_$1I4152_wr_clk , _6I4412_$1I4152_rd_en , _6I4412_$1I4152_rd_clk , _6I4412_$1I4152_ainit , _6I4412_$1I4152_dout , _6I4412_$1I4152_full , _6I4412_$1I4152_empty  );

// ----------------------------------- //

 wire  _6I4412_$1I3863_CHBONDDONE;

 wire [3:0] _6I4412_$1I3863_CHBONDO;

 wire  _6I4412_$1I3863_CONFIGOUT;

 wire [1:0] _6I4412_$1I3863_RXBUFSTATUS;

 wire [3:0] _6I4412_$1I3863_RXCHARISCOMMA;

 wire [3:0] _6I4412_$1I3863_RXCHARISK;

 wire  _6I4412_$1I3863_RXCHECKINGCRC;

 wire [2:0] _6I4412_$1I3863_RXCLKCORCNT;

 wire  _6I4412_$1I3863_RXCOMMADET;

 wire  _6I4412_$1I3863_RXCRCERR;

 wire [31:0] _6I4412_$1I3863_RXDATA;

 wire [3:0] _6I4412_$1I3863_RXDISPERR;

 wire [1:0] _6I4412_$1I3863_RXLOSSOFSYNC;

 wire [3:0] _6I4412_$1I3863_RXNOTINTABLE;

 wire  _6I4412_$1I3863_RXREALIGN;

 wire  _6I4412_$1I3863_RXRECCLK;

 wire [3:0] _6I4412_$1I3863_RXRUNDISP;

 wire  _6I4412_$1I3863_TXBUFERR;

 wire [3:0] _6I4412_$1I3863_TXKERR;

 wire  _6I4412_$1I3863_TXN;

 wire  _6I4412_$1I3863_TXP;

 wire [3:0] _6I4412_$1I3863_TXRUNDISP;

 wire  _6I4412_$1I3863_BREFCLK;
 reg [1:16] _6I4412_$1I3863_BREFCLK__vlIN;
 cstw cstw_639 (_6I4412_$1I3863_BREFCLK, _6I4412_$1I3863_BREFCLK__vlIN);

 wire  _6I4412_$1I3863_BREFCLK2;
 reg [1:16] _6I4412_$1I3863_BREFCLK2__vlIN;
 cstw cstw_640 (_6I4412_$1I3863_BREFCLK2, _6I4412_$1I3863_BREFCLK2__vlIN);

 wire [3:0] _6I4412_$1I3863_CHBONDI;
 reg [1:16] _6I4412_$1I3863_CHBONDI_3__vlIN;
 cstw cstw_641_3 (_6I4412_$1I3863_CHBONDI[3], _6I4412_$1I3863_CHBONDI_3__vlIN);
 reg [1:16] _6I4412_$1I3863_CHBONDI_2__vlIN;
 cstw cstw_641_2 (_6I4412_$1I3863_CHBONDI[2], _6I4412_$1I3863_CHBONDI_2__vlIN);
 reg [1:16] _6I4412_$1I3863_CHBONDI_1__vlIN;
 cstw cstw_641_1 (_6I4412_$1I3863_CHBONDI[1], _6I4412_$1I3863_CHBONDI_1__vlIN);
 reg [1:16] _6I4412_$1I3863_CHBONDI_0__vlIN;
 cstw cstw_641_0 (_6I4412_$1I3863_CHBONDI[0], _6I4412_$1I3863_CHBONDI_0__vlIN);

 wire  _6I4412_$1I3863_CONFIGENABLE;
 reg [1:16] _6I4412_$1I3863_CONFIGENABLE__vlIN;
 cstw cstw_642 (_6I4412_$1I3863_CONFIGENABLE, _6I4412_$1I3863_CONFIGENABLE__vlIN);

 wire  _6I4412_$1I3863_CONFIGIN;
 reg [1:16] _6I4412_$1I3863_CONFIGIN__vlIN;
 cstw cstw_643 (_6I4412_$1I3863_CONFIGIN, _6I4412_$1I3863_CONFIGIN__vlIN);

 wire  _6I4412_$1I3863_ENCHANSYNC;
 reg [1:16] _6I4412_$1I3863_ENCHANSYNC__vlIN;
 cstw cstw_644 (_6I4412_$1I3863_ENCHANSYNC, _6I4412_$1I3863_ENCHANSYNC__vlIN);

 wire  _6I4412_$1I3863_ENMCOMMAALIGN;
 reg [1:16] _6I4412_$1I3863_ENMCOMMAALIGN__vlIN;
 cstw cstw_645 (_6I4412_$1I3863_ENMCOMMAALIGN, _6I4412_$1I3863_ENMCOMMAALIGN__vlIN);

 wire  _6I4412_$1I3863_ENPCOMMAALIGN;
 reg [1:16] _6I4412_$1I3863_ENPCOMMAALIGN__vlIN;
 cstw cstw_646 (_6I4412_$1I3863_ENPCOMMAALIGN, _6I4412_$1I3863_ENPCOMMAALIGN__vlIN);

 wire [1:0] _6I4412_$1I3863_LOOPBACK;
 reg [1:16] _6I4412_$1I3863_LOOPBACK_1__vlIN;
 cstw cstw_647_1 (_6I4412_$1I3863_LOOPBACK[1], _6I4412_$1I3863_LOOPBACK_1__vlIN);
 reg [1:16] _6I4412_$1I3863_LOOPBACK_0__vlIN;
 cstw cstw_647_0 (_6I4412_$1I3863_LOOPBACK[0], _6I4412_$1I3863_LOOPBACK_0__vlIN);

 wire  _6I4412_$1I3863_POWERDOWN;
 reg [1:16] _6I4412_$1I3863_POWERDOWN__vlIN;
 cstw cstw_648 (_6I4412_$1I3863_POWERDOWN, _6I4412_$1I3863_POWERDOWN__vlIN);

 wire  _6I4412_$1I3863_REFCLK;
 reg [1:16] _6I4412_$1I3863_REFCLK__vlIN;
 cstw cstw_649 (_6I4412_$1I3863_REFCLK, _6I4412_$1I3863_REFCLK__vlIN);

 wire  _6I4412_$1I3863_REFCLK2;
 reg [1:16] _6I4412_$1I3863_REFCLK2__vlIN;
 cstw cstw_650 (_6I4412_$1I3863_REFCLK2, _6I4412_$1I3863_REFCLK2__vlIN);

 wire  _6I4412_$1I3863_REFCLKSEL;
 reg [1:16] _6I4412_$1I3863_REFCLKSEL__vlIN;
 cstw cstw_651 (_6I4412_$1I3863_REFCLKSEL, _6I4412_$1I3863_REFCLKSEL__vlIN);

 wire  _6I4412_$1I3863_RXN;
 reg [1:16] _6I4412_$1I3863_RXN__vlIN;
 cstw cstw_652 (_6I4412_$1I3863_RXN, _6I4412_$1I3863_RXN__vlIN);

 wire  _6I4412_$1I3863_RXP;
 reg [1:16] _6I4412_$1I3863_RXP__vlIN;
 cstw cstw_653 (_6I4412_$1I3863_RXP, _6I4412_$1I3863_RXP__vlIN);

 wire  _6I4412_$1I3863_RXPOLARITY;
 reg [1:16] _6I4412_$1I3863_RXPOLARITY__vlIN;
 cstw cstw_654 (_6I4412_$1I3863_RXPOLARITY, _6I4412_$1I3863_RXPOLARITY__vlIN);

 wire  _6I4412_$1I3863_RXRESET;
 reg [1:16] _6I4412_$1I3863_RXRESET__vlIN;
 cstw cstw_655 (_6I4412_$1I3863_RXRESET, _6I4412_$1I3863_RXRESET__vlIN);

 wire  _6I4412_$1I3863_RXUSRCLK;
 reg [1:16] _6I4412_$1I3863_RXUSRCLK__vlIN;
 cstw cstw_656 (_6I4412_$1I3863_RXUSRCLK, _6I4412_$1I3863_RXUSRCLK__vlIN);

 wire  _6I4412_$1I3863_RXUSRCLK2;
 reg [1:16] _6I4412_$1I3863_RXUSRCLK2__vlIN;
 cstw cstw_657 (_6I4412_$1I3863_RXUSRCLK2, _6I4412_$1I3863_RXUSRCLK2__vlIN);

 wire [3:0] _6I4412_$1I3863_TXBYPASS8B10B;
 reg [1:16] _6I4412_$1I3863_TXBYPASS8B10B_3__vlIN;
 cstw cstw_658_3 (_6I4412_$1I3863_TXBYPASS8B10B[3], _6I4412_$1I3863_TXBYPASS8B10B_3__vlIN);
 reg [1:16] _6I4412_$1I3863_TXBYPASS8B10B_2__vlIN;
 cstw cstw_658_2 (_6I4412_$1I3863_TXBYPASS8B10B[2], _6I4412_$1I3863_TXBYPASS8B10B_2__vlIN);
 reg [1:16] _6I4412_$1I3863_TXBYPASS8B10B_1__vlIN;
 cstw cstw_658_1 (_6I4412_$1I3863_TXBYPASS8B10B[1], _6I4412_$1I3863_TXBYPASS8B10B_1__vlIN);
 reg [1:16] _6I4412_$1I3863_TXBYPASS8B10B_0__vlIN;
 cstw cstw_658_0 (_6I4412_$1I3863_TXBYPASS8B10B[0], _6I4412_$1I3863_TXBYPASS8B10B_0__vlIN);

 wire [3:0] _6I4412_$1I3863_TXCHARDISPMODE;
 reg [1:16] _6I4412_$1I3863_TXCHARDISPMODE_3__vlIN;
 cstw cstw_659_3 (_6I4412_$1I3863_TXCHARDISPMODE[3], _6I4412_$1I3863_TXCHARDISPMODE_3__vlIN);
 reg [1:16] _6I4412_$1I3863_TXCHARDISPMODE_2__vlIN;
 cstw cstw_659_2 (_6I4412_$1I3863_TXCHARDISPMODE[2], _6I4412_$1I3863_TXCHARDISPMODE_2__vlIN);
 reg [1:16] _6I4412_$1I3863_TXCHARDISPMODE_1__vlIN;
 cstw cstw_659_1 (_6I4412_$1I3863_TXCHARDISPMODE[1], _6I4412_$1I3863_TXCHARDISPMODE_1__vlIN);
 reg [1:16] _6I4412_$1I3863_TXCHARDISPMODE_0__vlIN;
 cstw cstw_659_0 (_6I4412_$1I3863_TXCHARDISPMODE[0], _6I4412_$1I3863_TXCHARDISPMODE_0__vlIN);

 wire [3:0] _6I4412_$1I3863_TXCHARDISPVAL;
 reg [1:16] _6I4412_$1I3863_TXCHARDISPVAL_3__vlIN;
 cstw cstw_660_3 (_6I4412_$1I3863_TXCHARDISPVAL[3], _6I4412_$1I3863_TXCHARDISPVAL_3__vlIN);
 reg [1:16] _6I4412_$1I3863_TXCHARDISPVAL_2__vlIN;
 cstw cstw_660_2 (_6I4412_$1I3863_TXCHARDISPVAL[2], _6I4412_$1I3863_TXCHARDISPVAL_2__vlIN);
 reg [1:16] _6I4412_$1I3863_TXCHARDISPVAL_1__vlIN;
 cstw cstw_660_1 (_6I4412_$1I3863_TXCHARDISPVAL[1], _6I4412_$1I3863_TXCHARDISPVAL_1__vlIN);
 reg [1:16] _6I4412_$1I3863_TXCHARDISPVAL_0__vlIN;
 cstw cstw_660_0 (_6I4412_$1I3863_TXCHARDISPVAL[0], _6I4412_$1I3863_TXCHARDISPVAL_0__vlIN);

 wire [3:0] _6I4412_$1I3863_TXCHARISK;
 reg [1:16] _6I4412_$1I3863_TXCHARISK_3__vlIN;
 cstw cstw_661_3 (_6I4412_$1I3863_TXCHARISK[3], _6I4412_$1I3863_TXCHARISK_3__vlIN);
 reg [1:16] _6I4412_$1I3863_TXCHARISK_2__vlIN;
 cstw cstw_661_2 (_6I4412_$1I3863_TXCHARISK[2], _6I4412_$1I3863_TXCHARISK_2__vlIN);
 reg [1:16] _6I4412_$1I3863_TXCHARISK_1__vlIN;
 cstw cstw_661_1 (_6I4412_$1I3863_TXCHARISK[1], _6I4412_$1I3863_TXCHARISK_1__vlIN);
 reg [1:16] _6I4412_$1I3863_TXCHARISK_0__vlIN;
 cstw cstw_661_0 (_6I4412_$1I3863_TXCHARISK[0], _6I4412_$1I3863_TXCHARISK_0__vlIN);

 wire [31:0] _6I4412_$1I3863_TXDATA;
 reg [1:16] _6I4412_$1I3863_TXDATA_31__vlIN;
 cstw cstw_662_31 (_6I4412_$1I3863_TXDATA[31], _6I4412_$1I3863_TXDATA_31__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_30__vlIN;
 cstw cstw_662_30 (_6I4412_$1I3863_TXDATA[30], _6I4412_$1I3863_TXDATA_30__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_29__vlIN;
 cstw cstw_662_29 (_6I4412_$1I3863_TXDATA[29], _6I4412_$1I3863_TXDATA_29__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_28__vlIN;
 cstw cstw_662_28 (_6I4412_$1I3863_TXDATA[28], _6I4412_$1I3863_TXDATA_28__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_27__vlIN;
 cstw cstw_662_27 (_6I4412_$1I3863_TXDATA[27], _6I4412_$1I3863_TXDATA_27__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_26__vlIN;
 cstw cstw_662_26 (_6I4412_$1I3863_TXDATA[26], _6I4412_$1I3863_TXDATA_26__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_25__vlIN;
 cstw cstw_662_25 (_6I4412_$1I3863_TXDATA[25], _6I4412_$1I3863_TXDATA_25__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_24__vlIN;
 cstw cstw_662_24 (_6I4412_$1I3863_TXDATA[24], _6I4412_$1I3863_TXDATA_24__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_23__vlIN;
 cstw cstw_662_23 (_6I4412_$1I3863_TXDATA[23], _6I4412_$1I3863_TXDATA_23__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_22__vlIN;
 cstw cstw_662_22 (_6I4412_$1I3863_TXDATA[22], _6I4412_$1I3863_TXDATA_22__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_21__vlIN;
 cstw cstw_662_21 (_6I4412_$1I3863_TXDATA[21], _6I4412_$1I3863_TXDATA_21__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_20__vlIN;
 cstw cstw_662_20 (_6I4412_$1I3863_TXDATA[20], _6I4412_$1I3863_TXDATA_20__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_19__vlIN;
 cstw cstw_662_19 (_6I4412_$1I3863_TXDATA[19], _6I4412_$1I3863_TXDATA_19__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_18__vlIN;
 cstw cstw_662_18 (_6I4412_$1I3863_TXDATA[18], _6I4412_$1I3863_TXDATA_18__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_17__vlIN;
 cstw cstw_662_17 (_6I4412_$1I3863_TXDATA[17], _6I4412_$1I3863_TXDATA_17__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_16__vlIN;
 cstw cstw_662_16 (_6I4412_$1I3863_TXDATA[16], _6I4412_$1I3863_TXDATA_16__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_15__vlIN;
 cstw cstw_662_15 (_6I4412_$1I3863_TXDATA[15], _6I4412_$1I3863_TXDATA_15__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_14__vlIN;
 cstw cstw_662_14 (_6I4412_$1I3863_TXDATA[14], _6I4412_$1I3863_TXDATA_14__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_13__vlIN;
 cstw cstw_662_13 (_6I4412_$1I3863_TXDATA[13], _6I4412_$1I3863_TXDATA_13__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_12__vlIN;
 cstw cstw_662_12 (_6I4412_$1I3863_TXDATA[12], _6I4412_$1I3863_TXDATA_12__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_11__vlIN;
 cstw cstw_662_11 (_6I4412_$1I3863_TXDATA[11], _6I4412_$1I3863_TXDATA_11__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_10__vlIN;
 cstw cstw_662_10 (_6I4412_$1I3863_TXDATA[10], _6I4412_$1I3863_TXDATA_10__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_9__vlIN;
 cstw cstw_662_9 (_6I4412_$1I3863_TXDATA[9], _6I4412_$1I3863_TXDATA_9__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_8__vlIN;
 cstw cstw_662_8 (_6I4412_$1I3863_TXDATA[8], _6I4412_$1I3863_TXDATA_8__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_7__vlIN;
 cstw cstw_662_7 (_6I4412_$1I3863_TXDATA[7], _6I4412_$1I3863_TXDATA_7__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_6__vlIN;
 cstw cstw_662_6 (_6I4412_$1I3863_TXDATA[6], _6I4412_$1I3863_TXDATA_6__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_5__vlIN;
 cstw cstw_662_5 (_6I4412_$1I3863_TXDATA[5], _6I4412_$1I3863_TXDATA_5__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_4__vlIN;
 cstw cstw_662_4 (_6I4412_$1I3863_TXDATA[4], _6I4412_$1I3863_TXDATA_4__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_3__vlIN;
 cstw cstw_662_3 (_6I4412_$1I3863_TXDATA[3], _6I4412_$1I3863_TXDATA_3__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_2__vlIN;
 cstw cstw_662_2 (_6I4412_$1I3863_TXDATA[2], _6I4412_$1I3863_TXDATA_2__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_1__vlIN;
 cstw cstw_662_1 (_6I4412_$1I3863_TXDATA[1], _6I4412_$1I3863_TXDATA_1__vlIN);
 reg [1:16] _6I4412_$1I3863_TXDATA_0__vlIN;
 cstw cstw_662_0 (_6I4412_$1I3863_TXDATA[0], _6I4412_$1I3863_TXDATA_0__vlIN);

 wire  _6I4412_$1I3863_TXFORCECRCERR;
 reg [1:16] _6I4412_$1I3863_TXFORCECRCERR__vlIN;
 cstw cstw_663 (_6I4412_$1I3863_TXFORCECRCERR, _6I4412_$1I3863_TXFORCECRCERR__vlIN);

 wire  _6I4412_$1I3863_TXINHIBIT;
 reg [1:16] _6I4412_$1I3863_TXINHIBIT__vlIN;
 cstw cstw_664 (_6I4412_$1I3863_TXINHIBIT, _6I4412_$1I3863_TXINHIBIT__vlIN);

 wire  _6I4412_$1I3863_TXPOLARITY;
 reg [1:16] _6I4412_$1I3863_TXPOLARITY__vlIN;
 cstw cstw_665 (_6I4412_$1I3863_TXPOLARITY, _6I4412_$1I3863_TXPOLARITY__vlIN);

 wire  _6I4412_$1I3863_TXRESET;
 reg [1:16] _6I4412_$1I3863_TXRESET__vlIN;
 cstw cstw_666 (_6I4412_$1I3863_TXRESET, _6I4412_$1I3863_TXRESET__vlIN);

 wire  _6I4412_$1I3863_TXUSRCLK;
 reg [1:16] _6I4412_$1I3863_TXUSRCLK__vlIN;
 cstw cstw_667 (_6I4412_$1I3863_TXUSRCLK, _6I4412_$1I3863_TXUSRCLK__vlIN);

 wire  _6I4412_$1I3863_TXUSRCLK2;
 reg [1:16] _6I4412_$1I3863_TXUSRCLK2__vlIN;
 cstw cstw_668 (_6I4412_$1I3863_TXUSRCLK2, _6I4412_$1I3863_TXUSRCLK2__vlIN);

 GT_CUSTOM _6I4412_$1I3863 ( _6I4412_$1I3863_CHBONDDONE , _6I4412_$1I3863_CHBONDO , _6I4412_$1I3863_CONFIGOUT , _6I4412_$1I3863_RXBUFSTATUS , _6I4412_$1I3863_RXCHARISCOMMA , _6I4412_$1I3863_RXCHARISK , _6I4412_$1I3863_RXCHECKINGCRC , _6I4412_$1I3863_RXCLKCORCNT , _6I4412_$1I3863_RXCOMMADET , _6I4412_$1I3863_RXCRCERR , _6I4412_$1I3863_RXDATA , _6I4412_$1I3863_RXDISPERR , _6I4412_$1I3863_RXLOSSOFSYNC , _6I4412_$1I3863_RXNOTINTABLE , _6I4412_$1I3863_RXREALIGN , _6I4412_$1I3863_RXRECCLK , _6I4412_$1I3863_RXRUNDISP , _6I4412_$1I3863_TXBUFERR , _6I4412_$1I3863_TXKERR , _6I4412_$1I3863_TXN , _6I4412_$1I3863_TXP , _6I4412_$1I3863_TXRUNDISP , _6I4412_$1I3863_BREFCLK , _6I4412_$1I3863_BREFCLK2 , _6I4412_$1I3863_CHBONDI , _6I4412_$1I3863_CONFIGENABLE , _6I4412_$1I3863_CONFIGIN , _6I4412_$1I3863_ENCHANSYNC , _6I4412_$1I3863_ENMCOMMAALIGN , _6I4412_$1I3863_ENPCOMMAALIGN , _6I4412_$1I3863_LOOPBACK , _6I4412_$1I3863_POWERDOWN , _6I4412_$1I3863_REFCLK , _6I4412_$1I3863_REFCLK2 , _6I4412_$1I3863_REFCLKSEL , _6I4412_$1I3863_RXN , _6I4412_$1I3863_RXP , _6I4412_$1I3863_RXPOLARITY , _6I4412_$1I3863_RXRESET , _6I4412_$1I3863_RXUSRCLK , _6I4412_$1I3863_RXUSRCLK2 , _6I4412_$1I3863_TXBYPASS8B10B , _6I4412_$1I3863_TXCHARDISPMODE , _6I4412_$1I3863_TXCHARDISPVAL , _6I4412_$1I3863_TXCHARISK , _6I4412_$1I3863_TXDATA , _6I4412_$1I3863_TXFORCECRCERR , _6I4412_$1I3863_TXINHIBIT , _6I4412_$1I3863_TXPOLARITY , _6I4412_$1I3863_TXRESET , _6I4412_$1I3863_TXUSRCLK , _6I4412_$1I3863_TXUSRCLK2  );

// ----------------------------------- //

 wire [7:0] _6I4143_$1I4488_$1I4621_DOA;

 wire [15:0] _6I4143_$1I4488_$1I4621_DOB;

 wire [0:0] _6I4143_$1I4488_$1I4621_DOPA;

 wire [1:0] _6I4143_$1I4488_$1I4621_DOPB;

 wire [10:0] _6I4143_$1I4488_$1I4621_ADDRA;
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_669_10 (_6I4143_$1I4488_$1I4621_ADDRA[10], _6I4143_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_669_9 (_6I4143_$1I4488_$1I4621_ADDRA[9], _6I4143_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_669_8 (_6I4143_$1I4488_$1I4621_ADDRA[8], _6I4143_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_669_7 (_6I4143_$1I4488_$1I4621_ADDRA[7], _6I4143_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_669_6 (_6I4143_$1I4488_$1I4621_ADDRA[6], _6I4143_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_669_5 (_6I4143_$1I4488_$1I4621_ADDRA[5], _6I4143_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_669_4 (_6I4143_$1I4488_$1I4621_ADDRA[4], _6I4143_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_669_3 (_6I4143_$1I4488_$1I4621_ADDRA[3], _6I4143_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_669_2 (_6I4143_$1I4488_$1I4621_ADDRA[2], _6I4143_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_669_1 (_6I4143_$1I4488_$1I4621_ADDRA[1], _6I4143_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_669_0 (_6I4143_$1I4488_$1I4621_ADDRA[0], _6I4143_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _6I4143_$1I4488_$1I4621_ADDRB;
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_670_9 (_6I4143_$1I4488_$1I4621_ADDRB[9], _6I4143_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_670_8 (_6I4143_$1I4488_$1I4621_ADDRB[8], _6I4143_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_670_7 (_6I4143_$1I4488_$1I4621_ADDRB[7], _6I4143_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_670_6 (_6I4143_$1I4488_$1I4621_ADDRB[6], _6I4143_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_670_5 (_6I4143_$1I4488_$1I4621_ADDRB[5], _6I4143_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_670_4 (_6I4143_$1I4488_$1I4621_ADDRB[4], _6I4143_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_670_3 (_6I4143_$1I4488_$1I4621_ADDRB[3], _6I4143_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_670_2 (_6I4143_$1I4488_$1I4621_ADDRB[2], _6I4143_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_670_1 (_6I4143_$1I4488_$1I4621_ADDRB[1], _6I4143_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_670_0 (_6I4143_$1I4488_$1I4621_ADDRB[0], _6I4143_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _6I4143_$1I4488_$1I4621_CLKA;
 reg [1:16] _6I4143_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_671 (_6I4143_$1I4488_$1I4621_CLKA, _6I4143_$1I4488_$1I4621_CLKA__vlIN);

 wire  _6I4143_$1I4488_$1I4621_CLKB;
 reg [1:16] _6I4143_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_672 (_6I4143_$1I4488_$1I4621_CLKB, _6I4143_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _6I4143_$1I4488_$1I4621_DIA;
 reg [1:16] _6I4143_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_673_7 (_6I4143_$1I4488_$1I4621_DIA[7], _6I4143_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_673_6 (_6I4143_$1I4488_$1I4621_DIA[6], _6I4143_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_673_5 (_6I4143_$1I4488_$1I4621_DIA[5], _6I4143_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_673_4 (_6I4143_$1I4488_$1I4621_DIA[4], _6I4143_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_673_3 (_6I4143_$1I4488_$1I4621_DIA[3], _6I4143_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_673_2 (_6I4143_$1I4488_$1I4621_DIA[2], _6I4143_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_673_1 (_6I4143_$1I4488_$1I4621_DIA[1], _6I4143_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_673_0 (_6I4143_$1I4488_$1I4621_DIA[0], _6I4143_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _6I4143_$1I4488_$1I4621_DIB;
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_674_15 (_6I4143_$1I4488_$1I4621_DIB[15], _6I4143_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_674_14 (_6I4143_$1I4488_$1I4621_DIB[14], _6I4143_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_674_13 (_6I4143_$1I4488_$1I4621_DIB[13], _6I4143_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_674_12 (_6I4143_$1I4488_$1I4621_DIB[12], _6I4143_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_674_11 (_6I4143_$1I4488_$1I4621_DIB[11], _6I4143_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_674_10 (_6I4143_$1I4488_$1I4621_DIB[10], _6I4143_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_674_9 (_6I4143_$1I4488_$1I4621_DIB[9], _6I4143_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_674_8 (_6I4143_$1I4488_$1I4621_DIB[8], _6I4143_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_674_7 (_6I4143_$1I4488_$1I4621_DIB[7], _6I4143_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_674_6 (_6I4143_$1I4488_$1I4621_DIB[6], _6I4143_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_674_5 (_6I4143_$1I4488_$1I4621_DIB[5], _6I4143_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_674_4 (_6I4143_$1I4488_$1I4621_DIB[4], _6I4143_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_674_3 (_6I4143_$1I4488_$1I4621_DIB[3], _6I4143_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_674_2 (_6I4143_$1I4488_$1I4621_DIB[2], _6I4143_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_674_1 (_6I4143_$1I4488_$1I4621_DIB[1], _6I4143_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_674_0 (_6I4143_$1I4488_$1I4621_DIB[0], _6I4143_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _6I4143_$1I4488_$1I4621_DIPA;
 reg [1:16] _6I4143_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_675_0 (_6I4143_$1I4488_$1I4621_DIPA[0], _6I4143_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _6I4143_$1I4488_$1I4621_DIPB;
 reg [1:16] _6I4143_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_676_1 (_6I4143_$1I4488_$1I4621_DIPB[1], _6I4143_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_676_0 (_6I4143_$1I4488_$1I4621_DIPB[0], _6I4143_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _6I4143_$1I4488_$1I4621_ENA;
 reg [1:16] _6I4143_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_677 (_6I4143_$1I4488_$1I4621_ENA, _6I4143_$1I4488_$1I4621_ENA__vlIN);

 wire  _6I4143_$1I4488_$1I4621_ENB;
 reg [1:16] _6I4143_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_678 (_6I4143_$1I4488_$1I4621_ENB, _6I4143_$1I4488_$1I4621_ENB__vlIN);

 wire  _6I4143_$1I4488_$1I4621_SSRA;
 reg [1:16] _6I4143_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_679 (_6I4143_$1I4488_$1I4621_SSRA, _6I4143_$1I4488_$1I4621_SSRA__vlIN);

 wire  _6I4143_$1I4488_$1I4621_SSRB;
 reg [1:16] _6I4143_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_680 (_6I4143_$1I4488_$1I4621_SSRB, _6I4143_$1I4488_$1I4621_SSRB__vlIN);

 wire  _6I4143_$1I4488_$1I4621_WEA;
 reg [1:16] _6I4143_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_681 (_6I4143_$1I4488_$1I4621_WEA, _6I4143_$1I4488_$1I4621_WEA__vlIN);

 wire  _6I4143_$1I4488_$1I4621_WEB;
 reg [1:16] _6I4143_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_682 (_6I4143_$1I4488_$1I4621_WEB, _6I4143_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _6I4143_$1I4488_$1I4621 ( _6I4143_$1I4488_$1I4621_DOA , _6I4143_$1I4488_$1I4621_DOB , _6I4143_$1I4488_$1I4621_DOPA , _6I4143_$1I4488_$1I4621_DOPB , _6I4143_$1I4488_$1I4621_ADDRA , _6I4143_$1I4488_$1I4621_ADDRB , _6I4143_$1I4488_$1I4621_CLKA , _6I4143_$1I4488_$1I4621_CLKB , _6I4143_$1I4488_$1I4621_DIA , _6I4143_$1I4488_$1I4621_DIB , _6I4143_$1I4488_$1I4621_DIPA , _6I4143_$1I4488_$1I4621_DIPB , _6I4143_$1I4488_$1I4621_ENA , _6I4143_$1I4488_$1I4621_ENB , _6I4143_$1I4488_$1I4621_SSRA , _6I4143_$1I4488_$1I4621_SSRB , _6I4143_$1I4488_$1I4621_WEA , _6I4143_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _6I4143_$1I4488_$1I4620_DOA;

 wire [15:0] _6I4143_$1I4488_$1I4620_DOB;

 wire [0:0] _6I4143_$1I4488_$1I4620_DOPA;

 wire [1:0] _6I4143_$1I4488_$1I4620_DOPB;

 wire [10:0] _6I4143_$1I4488_$1I4620_ADDRA;
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_683_10 (_6I4143_$1I4488_$1I4620_ADDRA[10], _6I4143_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_683_9 (_6I4143_$1I4488_$1I4620_ADDRA[9], _6I4143_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_683_8 (_6I4143_$1I4488_$1I4620_ADDRA[8], _6I4143_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_683_7 (_6I4143_$1I4488_$1I4620_ADDRA[7], _6I4143_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_683_6 (_6I4143_$1I4488_$1I4620_ADDRA[6], _6I4143_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_683_5 (_6I4143_$1I4488_$1I4620_ADDRA[5], _6I4143_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_683_4 (_6I4143_$1I4488_$1I4620_ADDRA[4], _6I4143_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_683_3 (_6I4143_$1I4488_$1I4620_ADDRA[3], _6I4143_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_683_2 (_6I4143_$1I4488_$1I4620_ADDRA[2], _6I4143_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_683_1 (_6I4143_$1I4488_$1I4620_ADDRA[1], _6I4143_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_683_0 (_6I4143_$1I4488_$1I4620_ADDRA[0], _6I4143_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _6I4143_$1I4488_$1I4620_ADDRB;
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_684_9 (_6I4143_$1I4488_$1I4620_ADDRB[9], _6I4143_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_684_8 (_6I4143_$1I4488_$1I4620_ADDRB[8], _6I4143_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_684_7 (_6I4143_$1I4488_$1I4620_ADDRB[7], _6I4143_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_684_6 (_6I4143_$1I4488_$1I4620_ADDRB[6], _6I4143_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_684_5 (_6I4143_$1I4488_$1I4620_ADDRB[5], _6I4143_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_684_4 (_6I4143_$1I4488_$1I4620_ADDRB[4], _6I4143_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_684_3 (_6I4143_$1I4488_$1I4620_ADDRB[3], _6I4143_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_684_2 (_6I4143_$1I4488_$1I4620_ADDRB[2], _6I4143_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_684_1 (_6I4143_$1I4488_$1I4620_ADDRB[1], _6I4143_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_684_0 (_6I4143_$1I4488_$1I4620_ADDRB[0], _6I4143_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _6I4143_$1I4488_$1I4620_CLKA;
 reg [1:16] _6I4143_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_685 (_6I4143_$1I4488_$1I4620_CLKA, _6I4143_$1I4488_$1I4620_CLKA__vlIN);

 wire  _6I4143_$1I4488_$1I4620_CLKB;
 reg [1:16] _6I4143_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_686 (_6I4143_$1I4488_$1I4620_CLKB, _6I4143_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _6I4143_$1I4488_$1I4620_DIA;
 reg [1:16] _6I4143_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_687_7 (_6I4143_$1I4488_$1I4620_DIA[7], _6I4143_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_687_6 (_6I4143_$1I4488_$1I4620_DIA[6], _6I4143_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_687_5 (_6I4143_$1I4488_$1I4620_DIA[5], _6I4143_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_687_4 (_6I4143_$1I4488_$1I4620_DIA[4], _6I4143_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_687_3 (_6I4143_$1I4488_$1I4620_DIA[3], _6I4143_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_687_2 (_6I4143_$1I4488_$1I4620_DIA[2], _6I4143_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_687_1 (_6I4143_$1I4488_$1I4620_DIA[1], _6I4143_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_687_0 (_6I4143_$1I4488_$1I4620_DIA[0], _6I4143_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _6I4143_$1I4488_$1I4620_DIB;
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_688_15 (_6I4143_$1I4488_$1I4620_DIB[15], _6I4143_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_688_14 (_6I4143_$1I4488_$1I4620_DIB[14], _6I4143_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_688_13 (_6I4143_$1I4488_$1I4620_DIB[13], _6I4143_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_688_12 (_6I4143_$1I4488_$1I4620_DIB[12], _6I4143_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_688_11 (_6I4143_$1I4488_$1I4620_DIB[11], _6I4143_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_688_10 (_6I4143_$1I4488_$1I4620_DIB[10], _6I4143_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_688_9 (_6I4143_$1I4488_$1I4620_DIB[9], _6I4143_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_688_8 (_6I4143_$1I4488_$1I4620_DIB[8], _6I4143_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_688_7 (_6I4143_$1I4488_$1I4620_DIB[7], _6I4143_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_688_6 (_6I4143_$1I4488_$1I4620_DIB[6], _6I4143_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_688_5 (_6I4143_$1I4488_$1I4620_DIB[5], _6I4143_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_688_4 (_6I4143_$1I4488_$1I4620_DIB[4], _6I4143_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_688_3 (_6I4143_$1I4488_$1I4620_DIB[3], _6I4143_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_688_2 (_6I4143_$1I4488_$1I4620_DIB[2], _6I4143_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_688_1 (_6I4143_$1I4488_$1I4620_DIB[1], _6I4143_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_688_0 (_6I4143_$1I4488_$1I4620_DIB[0], _6I4143_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _6I4143_$1I4488_$1I4620_DIPA;
 reg [1:16] _6I4143_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_689_0 (_6I4143_$1I4488_$1I4620_DIPA[0], _6I4143_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _6I4143_$1I4488_$1I4620_DIPB;
 reg [1:16] _6I4143_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_690_1 (_6I4143_$1I4488_$1I4620_DIPB[1], _6I4143_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _6I4143_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_690_0 (_6I4143_$1I4488_$1I4620_DIPB[0], _6I4143_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _6I4143_$1I4488_$1I4620_ENA;
 reg [1:16] _6I4143_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_691 (_6I4143_$1I4488_$1I4620_ENA, _6I4143_$1I4488_$1I4620_ENA__vlIN);

 wire  _6I4143_$1I4488_$1I4620_ENB;
 reg [1:16] _6I4143_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_692 (_6I4143_$1I4488_$1I4620_ENB, _6I4143_$1I4488_$1I4620_ENB__vlIN);

 wire  _6I4143_$1I4488_$1I4620_SSRA;
 reg [1:16] _6I4143_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_693 (_6I4143_$1I4488_$1I4620_SSRA, _6I4143_$1I4488_$1I4620_SSRA__vlIN);

 wire  _6I4143_$1I4488_$1I4620_SSRB;
 reg [1:16] _6I4143_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_694 (_6I4143_$1I4488_$1I4620_SSRB, _6I4143_$1I4488_$1I4620_SSRB__vlIN);

 wire  _6I4143_$1I4488_$1I4620_WEA;
 reg [1:16] _6I4143_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_695 (_6I4143_$1I4488_$1I4620_WEA, _6I4143_$1I4488_$1I4620_WEA__vlIN);

 wire  _6I4143_$1I4488_$1I4620_WEB;
 reg [1:16] _6I4143_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_696 (_6I4143_$1I4488_$1I4620_WEB, _6I4143_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _6I4143_$1I4488_$1I4620 ( _6I4143_$1I4488_$1I4620_DOA , _6I4143_$1I4488_$1I4620_DOB , _6I4143_$1I4488_$1I4620_DOPA , _6I4143_$1I4488_$1I4620_DOPB , _6I4143_$1I4488_$1I4620_ADDRA , _6I4143_$1I4488_$1I4620_ADDRB , _6I4143_$1I4488_$1I4620_CLKA , _6I4143_$1I4488_$1I4620_CLKB , _6I4143_$1I4488_$1I4620_DIA , _6I4143_$1I4488_$1I4620_DIB , _6I4143_$1I4488_$1I4620_DIPA , _6I4143_$1I4488_$1I4620_DIPB , _6I4143_$1I4488_$1I4620_ENA , _6I4143_$1I4488_$1I4620_ENB , _6I4143_$1I4488_$1I4620_SSRA , _6I4143_$1I4488_$1I4620_SSRB , _6I4143_$1I4488_$1I4620_WEA , _6I4143_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [4:0] _5I4382_$1I4152_din;
 reg [1:16] _5I4382_$1I4152_din_4__vlIN;
 cstw cstw_697_4 (_5I4382_$1I4152_din[4], _5I4382_$1I4152_din_4__vlIN);
 reg [1:16] _5I4382_$1I4152_din_3__vlIN;
 cstw cstw_697_3 (_5I4382_$1I4152_din[3], _5I4382_$1I4152_din_3__vlIN);
 reg [1:16] _5I4382_$1I4152_din_2__vlIN;
 cstw cstw_697_2 (_5I4382_$1I4152_din[2], _5I4382_$1I4152_din_2__vlIN);
 reg [1:16] _5I4382_$1I4152_din_1__vlIN;
 cstw cstw_697_1 (_5I4382_$1I4152_din[1], _5I4382_$1I4152_din_1__vlIN);
 reg [1:16] _5I4382_$1I4152_din_0__vlIN;
 cstw cstw_697_0 (_5I4382_$1I4152_din[0], _5I4382_$1I4152_din_0__vlIN);

 wire  _5I4382_$1I4152_wr_en;
 reg [1:16] _5I4382_$1I4152_wr_en__vlIN;
 cstw cstw_698 (_5I4382_$1I4152_wr_en, _5I4382_$1I4152_wr_en__vlIN);

 wire  _5I4382_$1I4152_wr_clk;
 reg [1:16] _5I4382_$1I4152_wr_clk__vlIN;
 cstw cstw_699 (_5I4382_$1I4152_wr_clk, _5I4382_$1I4152_wr_clk__vlIN);

 wire  _5I4382_$1I4152_rd_en;
 reg [1:16] _5I4382_$1I4152_rd_en__vlIN;
 cstw cstw_700 (_5I4382_$1I4152_rd_en, _5I4382_$1I4152_rd_en__vlIN);

 wire  _5I4382_$1I4152_rd_clk;
 reg [1:16] _5I4382_$1I4152_rd_clk__vlIN;
 cstw cstw_701 (_5I4382_$1I4152_rd_clk, _5I4382_$1I4152_rd_clk__vlIN);

 wire  _5I4382_$1I4152_ainit;
 reg [1:16] _5I4382_$1I4152_ainit__vlIN;
 cstw cstw_702 (_5I4382_$1I4152_ainit, _5I4382_$1I4152_ainit__vlIN);

 wire [4:0] _5I4382_$1I4152_dout;

 wire  _5I4382_$1I4152_full;

 wire  _5I4382_$1I4152_empty;

 af_clb_5x31rpm _5I4382_$1I4152 ( _5I4382_$1I4152_din , _5I4382_$1I4152_wr_en , _5I4382_$1I4152_wr_clk , _5I4382_$1I4152_rd_en , _5I4382_$1I4152_rd_clk , _5I4382_$1I4152_ainit , _5I4382_$1I4152_dout , _5I4382_$1I4152_full , _5I4382_$1I4152_empty  );

// ----------------------------------- //

 wire  _5I4382_$1I3863_CHBONDDONE;

 wire [3:0] _5I4382_$1I3863_CHBONDO;

 wire  _5I4382_$1I3863_CONFIGOUT;

 wire [1:0] _5I4382_$1I3863_RXBUFSTATUS;

 wire [3:0] _5I4382_$1I3863_RXCHARISCOMMA;

 wire [3:0] _5I4382_$1I3863_RXCHARISK;

 wire  _5I4382_$1I3863_RXCHECKINGCRC;

 wire [2:0] _5I4382_$1I3863_RXCLKCORCNT;

 wire  _5I4382_$1I3863_RXCOMMADET;

 wire  _5I4382_$1I3863_RXCRCERR;

 wire [31:0] _5I4382_$1I3863_RXDATA;

 wire [3:0] _5I4382_$1I3863_RXDISPERR;

 wire [1:0] _5I4382_$1I3863_RXLOSSOFSYNC;

 wire [3:0] _5I4382_$1I3863_RXNOTINTABLE;

 wire  _5I4382_$1I3863_RXREALIGN;

 wire  _5I4382_$1I3863_RXRECCLK;

 wire [3:0] _5I4382_$1I3863_RXRUNDISP;

 wire  _5I4382_$1I3863_TXBUFERR;

 wire [3:0] _5I4382_$1I3863_TXKERR;

 wire  _5I4382_$1I3863_TXN;

 wire  _5I4382_$1I3863_TXP;

 wire [3:0] _5I4382_$1I3863_TXRUNDISP;

 wire  _5I4382_$1I3863_BREFCLK;
 reg [1:16] _5I4382_$1I3863_BREFCLK__vlIN;
 cstw cstw_703 (_5I4382_$1I3863_BREFCLK, _5I4382_$1I3863_BREFCLK__vlIN);

 wire  _5I4382_$1I3863_BREFCLK2;
 reg [1:16] _5I4382_$1I3863_BREFCLK2__vlIN;
 cstw cstw_704 (_5I4382_$1I3863_BREFCLK2, _5I4382_$1I3863_BREFCLK2__vlIN);

 wire [3:0] _5I4382_$1I3863_CHBONDI;
 reg [1:16] _5I4382_$1I3863_CHBONDI_3__vlIN;
 cstw cstw_705_3 (_5I4382_$1I3863_CHBONDI[3], _5I4382_$1I3863_CHBONDI_3__vlIN);
 reg [1:16] _5I4382_$1I3863_CHBONDI_2__vlIN;
 cstw cstw_705_2 (_5I4382_$1I3863_CHBONDI[2], _5I4382_$1I3863_CHBONDI_2__vlIN);
 reg [1:16] _5I4382_$1I3863_CHBONDI_1__vlIN;
 cstw cstw_705_1 (_5I4382_$1I3863_CHBONDI[1], _5I4382_$1I3863_CHBONDI_1__vlIN);
 reg [1:16] _5I4382_$1I3863_CHBONDI_0__vlIN;
 cstw cstw_705_0 (_5I4382_$1I3863_CHBONDI[0], _5I4382_$1I3863_CHBONDI_0__vlIN);

 wire  _5I4382_$1I3863_CONFIGENABLE;
 reg [1:16] _5I4382_$1I3863_CONFIGENABLE__vlIN;
 cstw cstw_706 (_5I4382_$1I3863_CONFIGENABLE, _5I4382_$1I3863_CONFIGENABLE__vlIN);

 wire  _5I4382_$1I3863_CONFIGIN;
 reg [1:16] _5I4382_$1I3863_CONFIGIN__vlIN;
 cstw cstw_707 (_5I4382_$1I3863_CONFIGIN, _5I4382_$1I3863_CONFIGIN__vlIN);

 wire  _5I4382_$1I3863_ENCHANSYNC;
 reg [1:16] _5I4382_$1I3863_ENCHANSYNC__vlIN;
 cstw cstw_708 (_5I4382_$1I3863_ENCHANSYNC, _5I4382_$1I3863_ENCHANSYNC__vlIN);

 wire  _5I4382_$1I3863_ENMCOMMAALIGN;
 reg [1:16] _5I4382_$1I3863_ENMCOMMAALIGN__vlIN;
 cstw cstw_709 (_5I4382_$1I3863_ENMCOMMAALIGN, _5I4382_$1I3863_ENMCOMMAALIGN__vlIN);

 wire  _5I4382_$1I3863_ENPCOMMAALIGN;
 reg [1:16] _5I4382_$1I3863_ENPCOMMAALIGN__vlIN;
 cstw cstw_710 (_5I4382_$1I3863_ENPCOMMAALIGN, _5I4382_$1I3863_ENPCOMMAALIGN__vlIN);

 wire [1:0] _5I4382_$1I3863_LOOPBACK;
 reg [1:16] _5I4382_$1I3863_LOOPBACK_1__vlIN;
 cstw cstw_711_1 (_5I4382_$1I3863_LOOPBACK[1], _5I4382_$1I3863_LOOPBACK_1__vlIN);
 reg [1:16] _5I4382_$1I3863_LOOPBACK_0__vlIN;
 cstw cstw_711_0 (_5I4382_$1I3863_LOOPBACK[0], _5I4382_$1I3863_LOOPBACK_0__vlIN);

 wire  _5I4382_$1I3863_POWERDOWN;
 reg [1:16] _5I4382_$1I3863_POWERDOWN__vlIN;
 cstw cstw_712 (_5I4382_$1I3863_POWERDOWN, _5I4382_$1I3863_POWERDOWN__vlIN);

 wire  _5I4382_$1I3863_REFCLK;
 reg [1:16] _5I4382_$1I3863_REFCLK__vlIN;
 cstw cstw_713 (_5I4382_$1I3863_REFCLK, _5I4382_$1I3863_REFCLK__vlIN);

 wire  _5I4382_$1I3863_REFCLK2;
 reg [1:16] _5I4382_$1I3863_REFCLK2__vlIN;
 cstw cstw_714 (_5I4382_$1I3863_REFCLK2, _5I4382_$1I3863_REFCLK2__vlIN);

 wire  _5I4382_$1I3863_REFCLKSEL;
 reg [1:16] _5I4382_$1I3863_REFCLKSEL__vlIN;
 cstw cstw_715 (_5I4382_$1I3863_REFCLKSEL, _5I4382_$1I3863_REFCLKSEL__vlIN);

 wire  _5I4382_$1I3863_RXN;
 reg [1:16] _5I4382_$1I3863_RXN__vlIN;
 cstw cstw_716 (_5I4382_$1I3863_RXN, _5I4382_$1I3863_RXN__vlIN);

 wire  _5I4382_$1I3863_RXP;
 reg [1:16] _5I4382_$1I3863_RXP__vlIN;
 cstw cstw_717 (_5I4382_$1I3863_RXP, _5I4382_$1I3863_RXP__vlIN);

 wire  _5I4382_$1I3863_RXPOLARITY;
 reg [1:16] _5I4382_$1I3863_RXPOLARITY__vlIN;
 cstw cstw_718 (_5I4382_$1I3863_RXPOLARITY, _5I4382_$1I3863_RXPOLARITY__vlIN);

 wire  _5I4382_$1I3863_RXRESET;
 reg [1:16] _5I4382_$1I3863_RXRESET__vlIN;
 cstw cstw_719 (_5I4382_$1I3863_RXRESET, _5I4382_$1I3863_RXRESET__vlIN);

 wire  _5I4382_$1I3863_RXUSRCLK;
 reg [1:16] _5I4382_$1I3863_RXUSRCLK__vlIN;
 cstw cstw_720 (_5I4382_$1I3863_RXUSRCLK, _5I4382_$1I3863_RXUSRCLK__vlIN);

 wire  _5I4382_$1I3863_RXUSRCLK2;
 reg [1:16] _5I4382_$1I3863_RXUSRCLK2__vlIN;
 cstw cstw_721 (_5I4382_$1I3863_RXUSRCLK2, _5I4382_$1I3863_RXUSRCLK2__vlIN);

 wire [3:0] _5I4382_$1I3863_TXBYPASS8B10B;
 reg [1:16] _5I4382_$1I3863_TXBYPASS8B10B_3__vlIN;
 cstw cstw_722_3 (_5I4382_$1I3863_TXBYPASS8B10B[3], _5I4382_$1I3863_TXBYPASS8B10B_3__vlIN);
 reg [1:16] _5I4382_$1I3863_TXBYPASS8B10B_2__vlIN;
 cstw cstw_722_2 (_5I4382_$1I3863_TXBYPASS8B10B[2], _5I4382_$1I3863_TXBYPASS8B10B_2__vlIN);
 reg [1:16] _5I4382_$1I3863_TXBYPASS8B10B_1__vlIN;
 cstw cstw_722_1 (_5I4382_$1I3863_TXBYPASS8B10B[1], _5I4382_$1I3863_TXBYPASS8B10B_1__vlIN);
 reg [1:16] _5I4382_$1I3863_TXBYPASS8B10B_0__vlIN;
 cstw cstw_722_0 (_5I4382_$1I3863_TXBYPASS8B10B[0], _5I4382_$1I3863_TXBYPASS8B10B_0__vlIN);

 wire [3:0] _5I4382_$1I3863_TXCHARDISPMODE;
 reg [1:16] _5I4382_$1I3863_TXCHARDISPMODE_3__vlIN;
 cstw cstw_723_3 (_5I4382_$1I3863_TXCHARDISPMODE[3], _5I4382_$1I3863_TXCHARDISPMODE_3__vlIN);
 reg [1:16] _5I4382_$1I3863_TXCHARDISPMODE_2__vlIN;
 cstw cstw_723_2 (_5I4382_$1I3863_TXCHARDISPMODE[2], _5I4382_$1I3863_TXCHARDISPMODE_2__vlIN);
 reg [1:16] _5I4382_$1I3863_TXCHARDISPMODE_1__vlIN;
 cstw cstw_723_1 (_5I4382_$1I3863_TXCHARDISPMODE[1], _5I4382_$1I3863_TXCHARDISPMODE_1__vlIN);
 reg [1:16] _5I4382_$1I3863_TXCHARDISPMODE_0__vlIN;
 cstw cstw_723_0 (_5I4382_$1I3863_TXCHARDISPMODE[0], _5I4382_$1I3863_TXCHARDISPMODE_0__vlIN);

 wire [3:0] _5I4382_$1I3863_TXCHARDISPVAL;
 reg [1:16] _5I4382_$1I3863_TXCHARDISPVAL_3__vlIN;
 cstw cstw_724_3 (_5I4382_$1I3863_TXCHARDISPVAL[3], _5I4382_$1I3863_TXCHARDISPVAL_3__vlIN);
 reg [1:16] _5I4382_$1I3863_TXCHARDISPVAL_2__vlIN;
 cstw cstw_724_2 (_5I4382_$1I3863_TXCHARDISPVAL[2], _5I4382_$1I3863_TXCHARDISPVAL_2__vlIN);
 reg [1:16] _5I4382_$1I3863_TXCHARDISPVAL_1__vlIN;
 cstw cstw_724_1 (_5I4382_$1I3863_TXCHARDISPVAL[1], _5I4382_$1I3863_TXCHARDISPVAL_1__vlIN);
 reg [1:16] _5I4382_$1I3863_TXCHARDISPVAL_0__vlIN;
 cstw cstw_724_0 (_5I4382_$1I3863_TXCHARDISPVAL[0], _5I4382_$1I3863_TXCHARDISPVAL_0__vlIN);

 wire [3:0] _5I4382_$1I3863_TXCHARISK;
 reg [1:16] _5I4382_$1I3863_TXCHARISK_3__vlIN;
 cstw cstw_725_3 (_5I4382_$1I3863_TXCHARISK[3], _5I4382_$1I3863_TXCHARISK_3__vlIN);
 reg [1:16] _5I4382_$1I3863_TXCHARISK_2__vlIN;
 cstw cstw_725_2 (_5I4382_$1I3863_TXCHARISK[2], _5I4382_$1I3863_TXCHARISK_2__vlIN);
 reg [1:16] _5I4382_$1I3863_TXCHARISK_1__vlIN;
 cstw cstw_725_1 (_5I4382_$1I3863_TXCHARISK[1], _5I4382_$1I3863_TXCHARISK_1__vlIN);
 reg [1:16] _5I4382_$1I3863_TXCHARISK_0__vlIN;
 cstw cstw_725_0 (_5I4382_$1I3863_TXCHARISK[0], _5I4382_$1I3863_TXCHARISK_0__vlIN);

 wire [31:0] _5I4382_$1I3863_TXDATA;
 reg [1:16] _5I4382_$1I3863_TXDATA_31__vlIN;
 cstw cstw_726_31 (_5I4382_$1I3863_TXDATA[31], _5I4382_$1I3863_TXDATA_31__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_30__vlIN;
 cstw cstw_726_30 (_5I4382_$1I3863_TXDATA[30], _5I4382_$1I3863_TXDATA_30__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_29__vlIN;
 cstw cstw_726_29 (_5I4382_$1I3863_TXDATA[29], _5I4382_$1I3863_TXDATA_29__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_28__vlIN;
 cstw cstw_726_28 (_5I4382_$1I3863_TXDATA[28], _5I4382_$1I3863_TXDATA_28__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_27__vlIN;
 cstw cstw_726_27 (_5I4382_$1I3863_TXDATA[27], _5I4382_$1I3863_TXDATA_27__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_26__vlIN;
 cstw cstw_726_26 (_5I4382_$1I3863_TXDATA[26], _5I4382_$1I3863_TXDATA_26__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_25__vlIN;
 cstw cstw_726_25 (_5I4382_$1I3863_TXDATA[25], _5I4382_$1I3863_TXDATA_25__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_24__vlIN;
 cstw cstw_726_24 (_5I4382_$1I3863_TXDATA[24], _5I4382_$1I3863_TXDATA_24__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_23__vlIN;
 cstw cstw_726_23 (_5I4382_$1I3863_TXDATA[23], _5I4382_$1I3863_TXDATA_23__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_22__vlIN;
 cstw cstw_726_22 (_5I4382_$1I3863_TXDATA[22], _5I4382_$1I3863_TXDATA_22__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_21__vlIN;
 cstw cstw_726_21 (_5I4382_$1I3863_TXDATA[21], _5I4382_$1I3863_TXDATA_21__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_20__vlIN;
 cstw cstw_726_20 (_5I4382_$1I3863_TXDATA[20], _5I4382_$1I3863_TXDATA_20__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_19__vlIN;
 cstw cstw_726_19 (_5I4382_$1I3863_TXDATA[19], _5I4382_$1I3863_TXDATA_19__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_18__vlIN;
 cstw cstw_726_18 (_5I4382_$1I3863_TXDATA[18], _5I4382_$1I3863_TXDATA_18__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_17__vlIN;
 cstw cstw_726_17 (_5I4382_$1I3863_TXDATA[17], _5I4382_$1I3863_TXDATA_17__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_16__vlIN;
 cstw cstw_726_16 (_5I4382_$1I3863_TXDATA[16], _5I4382_$1I3863_TXDATA_16__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_15__vlIN;
 cstw cstw_726_15 (_5I4382_$1I3863_TXDATA[15], _5I4382_$1I3863_TXDATA_15__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_14__vlIN;
 cstw cstw_726_14 (_5I4382_$1I3863_TXDATA[14], _5I4382_$1I3863_TXDATA_14__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_13__vlIN;
 cstw cstw_726_13 (_5I4382_$1I3863_TXDATA[13], _5I4382_$1I3863_TXDATA_13__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_12__vlIN;
 cstw cstw_726_12 (_5I4382_$1I3863_TXDATA[12], _5I4382_$1I3863_TXDATA_12__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_11__vlIN;
 cstw cstw_726_11 (_5I4382_$1I3863_TXDATA[11], _5I4382_$1I3863_TXDATA_11__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_10__vlIN;
 cstw cstw_726_10 (_5I4382_$1I3863_TXDATA[10], _5I4382_$1I3863_TXDATA_10__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_9__vlIN;
 cstw cstw_726_9 (_5I4382_$1I3863_TXDATA[9], _5I4382_$1I3863_TXDATA_9__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_8__vlIN;
 cstw cstw_726_8 (_5I4382_$1I3863_TXDATA[8], _5I4382_$1I3863_TXDATA_8__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_7__vlIN;
 cstw cstw_726_7 (_5I4382_$1I3863_TXDATA[7], _5I4382_$1I3863_TXDATA_7__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_6__vlIN;
 cstw cstw_726_6 (_5I4382_$1I3863_TXDATA[6], _5I4382_$1I3863_TXDATA_6__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_5__vlIN;
 cstw cstw_726_5 (_5I4382_$1I3863_TXDATA[5], _5I4382_$1I3863_TXDATA_5__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_4__vlIN;
 cstw cstw_726_4 (_5I4382_$1I3863_TXDATA[4], _5I4382_$1I3863_TXDATA_4__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_3__vlIN;
 cstw cstw_726_3 (_5I4382_$1I3863_TXDATA[3], _5I4382_$1I3863_TXDATA_3__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_2__vlIN;
 cstw cstw_726_2 (_5I4382_$1I3863_TXDATA[2], _5I4382_$1I3863_TXDATA_2__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_1__vlIN;
 cstw cstw_726_1 (_5I4382_$1I3863_TXDATA[1], _5I4382_$1I3863_TXDATA_1__vlIN);
 reg [1:16] _5I4382_$1I3863_TXDATA_0__vlIN;
 cstw cstw_726_0 (_5I4382_$1I3863_TXDATA[0], _5I4382_$1I3863_TXDATA_0__vlIN);

 wire  _5I4382_$1I3863_TXFORCECRCERR;
 reg [1:16] _5I4382_$1I3863_TXFORCECRCERR__vlIN;
 cstw cstw_727 (_5I4382_$1I3863_TXFORCECRCERR, _5I4382_$1I3863_TXFORCECRCERR__vlIN);

 wire  _5I4382_$1I3863_TXINHIBIT;
 reg [1:16] _5I4382_$1I3863_TXINHIBIT__vlIN;
 cstw cstw_728 (_5I4382_$1I3863_TXINHIBIT, _5I4382_$1I3863_TXINHIBIT__vlIN);

 wire  _5I4382_$1I3863_TXPOLARITY;
 reg [1:16] _5I4382_$1I3863_TXPOLARITY__vlIN;
 cstw cstw_729 (_5I4382_$1I3863_TXPOLARITY, _5I4382_$1I3863_TXPOLARITY__vlIN);

 wire  _5I4382_$1I3863_TXRESET;
 reg [1:16] _5I4382_$1I3863_TXRESET__vlIN;
 cstw cstw_730 (_5I4382_$1I3863_TXRESET, _5I4382_$1I3863_TXRESET__vlIN);

 wire  _5I4382_$1I3863_TXUSRCLK;
 reg [1:16] _5I4382_$1I3863_TXUSRCLK__vlIN;
 cstw cstw_731 (_5I4382_$1I3863_TXUSRCLK, _5I4382_$1I3863_TXUSRCLK__vlIN);

 wire  _5I4382_$1I3863_TXUSRCLK2;
 reg [1:16] _5I4382_$1I3863_TXUSRCLK2__vlIN;
 cstw cstw_732 (_5I4382_$1I3863_TXUSRCLK2, _5I4382_$1I3863_TXUSRCLK2__vlIN);

 GT_CUSTOM _5I4382_$1I3863 ( _5I4382_$1I3863_CHBONDDONE , _5I4382_$1I3863_CHBONDO , _5I4382_$1I3863_CONFIGOUT , _5I4382_$1I3863_RXBUFSTATUS , _5I4382_$1I3863_RXCHARISCOMMA , _5I4382_$1I3863_RXCHARISK , _5I4382_$1I3863_RXCHECKINGCRC , _5I4382_$1I3863_RXCLKCORCNT , _5I4382_$1I3863_RXCOMMADET , _5I4382_$1I3863_RXCRCERR , _5I4382_$1I3863_RXDATA , _5I4382_$1I3863_RXDISPERR , _5I4382_$1I3863_RXLOSSOFSYNC , _5I4382_$1I3863_RXNOTINTABLE , _5I4382_$1I3863_RXREALIGN , _5I4382_$1I3863_RXRECCLK , _5I4382_$1I3863_RXRUNDISP , _5I4382_$1I3863_TXBUFERR , _5I4382_$1I3863_TXKERR , _5I4382_$1I3863_TXN , _5I4382_$1I3863_TXP , _5I4382_$1I3863_TXRUNDISP , _5I4382_$1I3863_BREFCLK , _5I4382_$1I3863_BREFCLK2 , _5I4382_$1I3863_CHBONDI , _5I4382_$1I3863_CONFIGENABLE , _5I4382_$1I3863_CONFIGIN , _5I4382_$1I3863_ENCHANSYNC , _5I4382_$1I3863_ENMCOMMAALIGN , _5I4382_$1I3863_ENPCOMMAALIGN , _5I4382_$1I3863_LOOPBACK , _5I4382_$1I3863_POWERDOWN , _5I4382_$1I3863_REFCLK , _5I4382_$1I3863_REFCLK2 , _5I4382_$1I3863_REFCLKSEL , _5I4382_$1I3863_RXN , _5I4382_$1I3863_RXP , _5I4382_$1I3863_RXPOLARITY , _5I4382_$1I3863_RXRESET , _5I4382_$1I3863_RXUSRCLK , _5I4382_$1I3863_RXUSRCLK2 , _5I4382_$1I3863_TXBYPASS8B10B , _5I4382_$1I3863_TXCHARDISPMODE , _5I4382_$1I3863_TXCHARDISPVAL , _5I4382_$1I3863_TXCHARISK , _5I4382_$1I3863_TXDATA , _5I4382_$1I3863_TXFORCECRCERR , _5I4382_$1I3863_TXINHIBIT , _5I4382_$1I3863_TXPOLARITY , _5I4382_$1I3863_TXRESET , _5I4382_$1I3863_TXUSRCLK , _5I4382_$1I3863_TXUSRCLK2  );

// ----------------------------------- //

 wire [7:0] _5I4143_$1I4488_$1I4621_DOA;

 wire [15:0] _5I4143_$1I4488_$1I4621_DOB;

 wire [0:0] _5I4143_$1I4488_$1I4621_DOPA;

 wire [1:0] _5I4143_$1I4488_$1I4621_DOPB;

 wire [10:0] _5I4143_$1I4488_$1I4621_ADDRA;
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_733_10 (_5I4143_$1I4488_$1I4621_ADDRA[10], _5I4143_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_733_9 (_5I4143_$1I4488_$1I4621_ADDRA[9], _5I4143_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_733_8 (_5I4143_$1I4488_$1I4621_ADDRA[8], _5I4143_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_733_7 (_5I4143_$1I4488_$1I4621_ADDRA[7], _5I4143_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_733_6 (_5I4143_$1I4488_$1I4621_ADDRA[6], _5I4143_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_733_5 (_5I4143_$1I4488_$1I4621_ADDRA[5], _5I4143_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_733_4 (_5I4143_$1I4488_$1I4621_ADDRA[4], _5I4143_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_733_3 (_5I4143_$1I4488_$1I4621_ADDRA[3], _5I4143_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_733_2 (_5I4143_$1I4488_$1I4621_ADDRA[2], _5I4143_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_733_1 (_5I4143_$1I4488_$1I4621_ADDRA[1], _5I4143_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_733_0 (_5I4143_$1I4488_$1I4621_ADDRA[0], _5I4143_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _5I4143_$1I4488_$1I4621_ADDRB;
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_734_9 (_5I4143_$1I4488_$1I4621_ADDRB[9], _5I4143_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_734_8 (_5I4143_$1I4488_$1I4621_ADDRB[8], _5I4143_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_734_7 (_5I4143_$1I4488_$1I4621_ADDRB[7], _5I4143_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_734_6 (_5I4143_$1I4488_$1I4621_ADDRB[6], _5I4143_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_734_5 (_5I4143_$1I4488_$1I4621_ADDRB[5], _5I4143_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_734_4 (_5I4143_$1I4488_$1I4621_ADDRB[4], _5I4143_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_734_3 (_5I4143_$1I4488_$1I4621_ADDRB[3], _5I4143_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_734_2 (_5I4143_$1I4488_$1I4621_ADDRB[2], _5I4143_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_734_1 (_5I4143_$1I4488_$1I4621_ADDRB[1], _5I4143_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_734_0 (_5I4143_$1I4488_$1I4621_ADDRB[0], _5I4143_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _5I4143_$1I4488_$1I4621_CLKA;
 reg [1:16] _5I4143_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_735 (_5I4143_$1I4488_$1I4621_CLKA, _5I4143_$1I4488_$1I4621_CLKA__vlIN);

 wire  _5I4143_$1I4488_$1I4621_CLKB;
 reg [1:16] _5I4143_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_736 (_5I4143_$1I4488_$1I4621_CLKB, _5I4143_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _5I4143_$1I4488_$1I4621_DIA;
 reg [1:16] _5I4143_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_737_7 (_5I4143_$1I4488_$1I4621_DIA[7], _5I4143_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_737_6 (_5I4143_$1I4488_$1I4621_DIA[6], _5I4143_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_737_5 (_5I4143_$1I4488_$1I4621_DIA[5], _5I4143_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_737_4 (_5I4143_$1I4488_$1I4621_DIA[4], _5I4143_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_737_3 (_5I4143_$1I4488_$1I4621_DIA[3], _5I4143_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_737_2 (_5I4143_$1I4488_$1I4621_DIA[2], _5I4143_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_737_1 (_5I4143_$1I4488_$1I4621_DIA[1], _5I4143_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_737_0 (_5I4143_$1I4488_$1I4621_DIA[0], _5I4143_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _5I4143_$1I4488_$1I4621_DIB;
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_738_15 (_5I4143_$1I4488_$1I4621_DIB[15], _5I4143_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_738_14 (_5I4143_$1I4488_$1I4621_DIB[14], _5I4143_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_738_13 (_5I4143_$1I4488_$1I4621_DIB[13], _5I4143_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_738_12 (_5I4143_$1I4488_$1I4621_DIB[12], _5I4143_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_738_11 (_5I4143_$1I4488_$1I4621_DIB[11], _5I4143_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_738_10 (_5I4143_$1I4488_$1I4621_DIB[10], _5I4143_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_738_9 (_5I4143_$1I4488_$1I4621_DIB[9], _5I4143_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_738_8 (_5I4143_$1I4488_$1I4621_DIB[8], _5I4143_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_738_7 (_5I4143_$1I4488_$1I4621_DIB[7], _5I4143_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_738_6 (_5I4143_$1I4488_$1I4621_DIB[6], _5I4143_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_738_5 (_5I4143_$1I4488_$1I4621_DIB[5], _5I4143_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_738_4 (_5I4143_$1I4488_$1I4621_DIB[4], _5I4143_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_738_3 (_5I4143_$1I4488_$1I4621_DIB[3], _5I4143_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_738_2 (_5I4143_$1I4488_$1I4621_DIB[2], _5I4143_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_738_1 (_5I4143_$1I4488_$1I4621_DIB[1], _5I4143_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_738_0 (_5I4143_$1I4488_$1I4621_DIB[0], _5I4143_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _5I4143_$1I4488_$1I4621_DIPA;
 reg [1:16] _5I4143_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_739_0 (_5I4143_$1I4488_$1I4621_DIPA[0], _5I4143_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _5I4143_$1I4488_$1I4621_DIPB;
 reg [1:16] _5I4143_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_740_1 (_5I4143_$1I4488_$1I4621_DIPB[1], _5I4143_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_740_0 (_5I4143_$1I4488_$1I4621_DIPB[0], _5I4143_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _5I4143_$1I4488_$1I4621_ENA;
 reg [1:16] _5I4143_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_741 (_5I4143_$1I4488_$1I4621_ENA, _5I4143_$1I4488_$1I4621_ENA__vlIN);

 wire  _5I4143_$1I4488_$1I4621_ENB;
 reg [1:16] _5I4143_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_742 (_5I4143_$1I4488_$1I4621_ENB, _5I4143_$1I4488_$1I4621_ENB__vlIN);

 wire  _5I4143_$1I4488_$1I4621_SSRA;
 reg [1:16] _5I4143_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_743 (_5I4143_$1I4488_$1I4621_SSRA, _5I4143_$1I4488_$1I4621_SSRA__vlIN);

 wire  _5I4143_$1I4488_$1I4621_SSRB;
 reg [1:16] _5I4143_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_744 (_5I4143_$1I4488_$1I4621_SSRB, _5I4143_$1I4488_$1I4621_SSRB__vlIN);

 wire  _5I4143_$1I4488_$1I4621_WEA;
 reg [1:16] _5I4143_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_745 (_5I4143_$1I4488_$1I4621_WEA, _5I4143_$1I4488_$1I4621_WEA__vlIN);

 wire  _5I4143_$1I4488_$1I4621_WEB;
 reg [1:16] _5I4143_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_746 (_5I4143_$1I4488_$1I4621_WEB, _5I4143_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _5I4143_$1I4488_$1I4621 ( _5I4143_$1I4488_$1I4621_DOA , _5I4143_$1I4488_$1I4621_DOB , _5I4143_$1I4488_$1I4621_DOPA , _5I4143_$1I4488_$1I4621_DOPB , _5I4143_$1I4488_$1I4621_ADDRA , _5I4143_$1I4488_$1I4621_ADDRB , _5I4143_$1I4488_$1I4621_CLKA , _5I4143_$1I4488_$1I4621_CLKB , _5I4143_$1I4488_$1I4621_DIA , _5I4143_$1I4488_$1I4621_DIB , _5I4143_$1I4488_$1I4621_DIPA , _5I4143_$1I4488_$1I4621_DIPB , _5I4143_$1I4488_$1I4621_ENA , _5I4143_$1I4488_$1I4621_ENB , _5I4143_$1I4488_$1I4621_SSRA , _5I4143_$1I4488_$1I4621_SSRB , _5I4143_$1I4488_$1I4621_WEA , _5I4143_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _5I4143_$1I4488_$1I4620_DOA;

 wire [15:0] _5I4143_$1I4488_$1I4620_DOB;

 wire [0:0] _5I4143_$1I4488_$1I4620_DOPA;

 wire [1:0] _5I4143_$1I4488_$1I4620_DOPB;

 wire [10:0] _5I4143_$1I4488_$1I4620_ADDRA;
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_747_10 (_5I4143_$1I4488_$1I4620_ADDRA[10], _5I4143_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_747_9 (_5I4143_$1I4488_$1I4620_ADDRA[9], _5I4143_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_747_8 (_5I4143_$1I4488_$1I4620_ADDRA[8], _5I4143_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_747_7 (_5I4143_$1I4488_$1I4620_ADDRA[7], _5I4143_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_747_6 (_5I4143_$1I4488_$1I4620_ADDRA[6], _5I4143_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_747_5 (_5I4143_$1I4488_$1I4620_ADDRA[5], _5I4143_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_747_4 (_5I4143_$1I4488_$1I4620_ADDRA[4], _5I4143_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_747_3 (_5I4143_$1I4488_$1I4620_ADDRA[3], _5I4143_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_747_2 (_5I4143_$1I4488_$1I4620_ADDRA[2], _5I4143_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_747_1 (_5I4143_$1I4488_$1I4620_ADDRA[1], _5I4143_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_747_0 (_5I4143_$1I4488_$1I4620_ADDRA[0], _5I4143_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _5I4143_$1I4488_$1I4620_ADDRB;
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_748_9 (_5I4143_$1I4488_$1I4620_ADDRB[9], _5I4143_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_748_8 (_5I4143_$1I4488_$1I4620_ADDRB[8], _5I4143_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_748_7 (_5I4143_$1I4488_$1I4620_ADDRB[7], _5I4143_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_748_6 (_5I4143_$1I4488_$1I4620_ADDRB[6], _5I4143_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_748_5 (_5I4143_$1I4488_$1I4620_ADDRB[5], _5I4143_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_748_4 (_5I4143_$1I4488_$1I4620_ADDRB[4], _5I4143_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_748_3 (_5I4143_$1I4488_$1I4620_ADDRB[3], _5I4143_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_748_2 (_5I4143_$1I4488_$1I4620_ADDRB[2], _5I4143_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_748_1 (_5I4143_$1I4488_$1I4620_ADDRB[1], _5I4143_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_748_0 (_5I4143_$1I4488_$1I4620_ADDRB[0], _5I4143_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _5I4143_$1I4488_$1I4620_CLKA;
 reg [1:16] _5I4143_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_749 (_5I4143_$1I4488_$1I4620_CLKA, _5I4143_$1I4488_$1I4620_CLKA__vlIN);

 wire  _5I4143_$1I4488_$1I4620_CLKB;
 reg [1:16] _5I4143_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_750 (_5I4143_$1I4488_$1I4620_CLKB, _5I4143_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _5I4143_$1I4488_$1I4620_DIA;
 reg [1:16] _5I4143_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_751_7 (_5I4143_$1I4488_$1I4620_DIA[7], _5I4143_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_751_6 (_5I4143_$1I4488_$1I4620_DIA[6], _5I4143_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_751_5 (_5I4143_$1I4488_$1I4620_DIA[5], _5I4143_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_751_4 (_5I4143_$1I4488_$1I4620_DIA[4], _5I4143_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_751_3 (_5I4143_$1I4488_$1I4620_DIA[3], _5I4143_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_751_2 (_5I4143_$1I4488_$1I4620_DIA[2], _5I4143_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_751_1 (_5I4143_$1I4488_$1I4620_DIA[1], _5I4143_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_751_0 (_5I4143_$1I4488_$1I4620_DIA[0], _5I4143_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _5I4143_$1I4488_$1I4620_DIB;
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_752_15 (_5I4143_$1I4488_$1I4620_DIB[15], _5I4143_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_752_14 (_5I4143_$1I4488_$1I4620_DIB[14], _5I4143_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_752_13 (_5I4143_$1I4488_$1I4620_DIB[13], _5I4143_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_752_12 (_5I4143_$1I4488_$1I4620_DIB[12], _5I4143_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_752_11 (_5I4143_$1I4488_$1I4620_DIB[11], _5I4143_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_752_10 (_5I4143_$1I4488_$1I4620_DIB[10], _5I4143_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_752_9 (_5I4143_$1I4488_$1I4620_DIB[9], _5I4143_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_752_8 (_5I4143_$1I4488_$1I4620_DIB[8], _5I4143_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_752_7 (_5I4143_$1I4488_$1I4620_DIB[7], _5I4143_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_752_6 (_5I4143_$1I4488_$1I4620_DIB[6], _5I4143_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_752_5 (_5I4143_$1I4488_$1I4620_DIB[5], _5I4143_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_752_4 (_5I4143_$1I4488_$1I4620_DIB[4], _5I4143_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_752_3 (_5I4143_$1I4488_$1I4620_DIB[3], _5I4143_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_752_2 (_5I4143_$1I4488_$1I4620_DIB[2], _5I4143_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_752_1 (_5I4143_$1I4488_$1I4620_DIB[1], _5I4143_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_752_0 (_5I4143_$1I4488_$1I4620_DIB[0], _5I4143_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _5I4143_$1I4488_$1I4620_DIPA;
 reg [1:16] _5I4143_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_753_0 (_5I4143_$1I4488_$1I4620_DIPA[0], _5I4143_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _5I4143_$1I4488_$1I4620_DIPB;
 reg [1:16] _5I4143_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_754_1 (_5I4143_$1I4488_$1I4620_DIPB[1], _5I4143_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _5I4143_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_754_0 (_5I4143_$1I4488_$1I4620_DIPB[0], _5I4143_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _5I4143_$1I4488_$1I4620_ENA;
 reg [1:16] _5I4143_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_755 (_5I4143_$1I4488_$1I4620_ENA, _5I4143_$1I4488_$1I4620_ENA__vlIN);

 wire  _5I4143_$1I4488_$1I4620_ENB;
 reg [1:16] _5I4143_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_756 (_5I4143_$1I4488_$1I4620_ENB, _5I4143_$1I4488_$1I4620_ENB__vlIN);

 wire  _5I4143_$1I4488_$1I4620_SSRA;
 reg [1:16] _5I4143_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_757 (_5I4143_$1I4488_$1I4620_SSRA, _5I4143_$1I4488_$1I4620_SSRA__vlIN);

 wire  _5I4143_$1I4488_$1I4620_SSRB;
 reg [1:16] _5I4143_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_758 (_5I4143_$1I4488_$1I4620_SSRB, _5I4143_$1I4488_$1I4620_SSRB__vlIN);

 wire  _5I4143_$1I4488_$1I4620_WEA;
 reg [1:16] _5I4143_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_759 (_5I4143_$1I4488_$1I4620_WEA, _5I4143_$1I4488_$1I4620_WEA__vlIN);

 wire  _5I4143_$1I4488_$1I4620_WEB;
 reg [1:16] _5I4143_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_760 (_5I4143_$1I4488_$1I4620_WEB, _5I4143_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _5I4143_$1I4488_$1I4620 ( _5I4143_$1I4488_$1I4620_DOA , _5I4143_$1I4488_$1I4620_DOB , _5I4143_$1I4488_$1I4620_DOPA , _5I4143_$1I4488_$1I4620_DOPB , _5I4143_$1I4488_$1I4620_ADDRA , _5I4143_$1I4488_$1I4620_ADDRB , _5I4143_$1I4488_$1I4620_CLKA , _5I4143_$1I4488_$1I4620_CLKB , _5I4143_$1I4488_$1I4620_DIA , _5I4143_$1I4488_$1I4620_DIB , _5I4143_$1I4488_$1I4620_DIPA , _5I4143_$1I4488_$1I4620_DIPB , _5I4143_$1I4488_$1I4620_ENA , _5I4143_$1I4488_$1I4620_ENB , _5I4143_$1I4488_$1I4620_SSRA , _5I4143_$1I4488_$1I4620_SSRB , _5I4143_$1I4488_$1I4620_WEA , _5I4143_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4657_$1I4488_$1I4621_DOA;

 wire [15:0] _4I4657_$1I4488_$1I4621_DOB;

 wire [0:0] _4I4657_$1I4488_$1I4621_DOPA;

 wire [1:0] _4I4657_$1I4488_$1I4621_DOPB;

 wire [10:0] _4I4657_$1I4488_$1I4621_ADDRA;
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_761_10 (_4I4657_$1I4488_$1I4621_ADDRA[10], _4I4657_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_761_9 (_4I4657_$1I4488_$1I4621_ADDRA[9], _4I4657_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_761_8 (_4I4657_$1I4488_$1I4621_ADDRA[8], _4I4657_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_761_7 (_4I4657_$1I4488_$1I4621_ADDRA[7], _4I4657_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_761_6 (_4I4657_$1I4488_$1I4621_ADDRA[6], _4I4657_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_761_5 (_4I4657_$1I4488_$1I4621_ADDRA[5], _4I4657_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_761_4 (_4I4657_$1I4488_$1I4621_ADDRA[4], _4I4657_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_761_3 (_4I4657_$1I4488_$1I4621_ADDRA[3], _4I4657_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_761_2 (_4I4657_$1I4488_$1I4621_ADDRA[2], _4I4657_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_761_1 (_4I4657_$1I4488_$1I4621_ADDRA[1], _4I4657_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_761_0 (_4I4657_$1I4488_$1I4621_ADDRA[0], _4I4657_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _4I4657_$1I4488_$1I4621_ADDRB;
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_762_9 (_4I4657_$1I4488_$1I4621_ADDRB[9], _4I4657_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_762_8 (_4I4657_$1I4488_$1I4621_ADDRB[8], _4I4657_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_762_7 (_4I4657_$1I4488_$1I4621_ADDRB[7], _4I4657_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_762_6 (_4I4657_$1I4488_$1I4621_ADDRB[6], _4I4657_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_762_5 (_4I4657_$1I4488_$1I4621_ADDRB[5], _4I4657_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_762_4 (_4I4657_$1I4488_$1I4621_ADDRB[4], _4I4657_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_762_3 (_4I4657_$1I4488_$1I4621_ADDRB[3], _4I4657_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_762_2 (_4I4657_$1I4488_$1I4621_ADDRB[2], _4I4657_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_762_1 (_4I4657_$1I4488_$1I4621_ADDRB[1], _4I4657_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_762_0 (_4I4657_$1I4488_$1I4621_ADDRB[0], _4I4657_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _4I4657_$1I4488_$1I4621_CLKA;
 reg [1:16] _4I4657_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_763 (_4I4657_$1I4488_$1I4621_CLKA, _4I4657_$1I4488_$1I4621_CLKA__vlIN);

 wire  _4I4657_$1I4488_$1I4621_CLKB;
 reg [1:16] _4I4657_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_764 (_4I4657_$1I4488_$1I4621_CLKB, _4I4657_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _4I4657_$1I4488_$1I4621_DIA;
 reg [1:16] _4I4657_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_765_7 (_4I4657_$1I4488_$1I4621_DIA[7], _4I4657_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_765_6 (_4I4657_$1I4488_$1I4621_DIA[6], _4I4657_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_765_5 (_4I4657_$1I4488_$1I4621_DIA[5], _4I4657_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_765_4 (_4I4657_$1I4488_$1I4621_DIA[4], _4I4657_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_765_3 (_4I4657_$1I4488_$1I4621_DIA[3], _4I4657_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_765_2 (_4I4657_$1I4488_$1I4621_DIA[2], _4I4657_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_765_1 (_4I4657_$1I4488_$1I4621_DIA[1], _4I4657_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_765_0 (_4I4657_$1I4488_$1I4621_DIA[0], _4I4657_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _4I4657_$1I4488_$1I4621_DIB;
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_766_15 (_4I4657_$1I4488_$1I4621_DIB[15], _4I4657_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_766_14 (_4I4657_$1I4488_$1I4621_DIB[14], _4I4657_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_766_13 (_4I4657_$1I4488_$1I4621_DIB[13], _4I4657_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_766_12 (_4I4657_$1I4488_$1I4621_DIB[12], _4I4657_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_766_11 (_4I4657_$1I4488_$1I4621_DIB[11], _4I4657_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_766_10 (_4I4657_$1I4488_$1I4621_DIB[10], _4I4657_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_766_9 (_4I4657_$1I4488_$1I4621_DIB[9], _4I4657_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_766_8 (_4I4657_$1I4488_$1I4621_DIB[8], _4I4657_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_766_7 (_4I4657_$1I4488_$1I4621_DIB[7], _4I4657_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_766_6 (_4I4657_$1I4488_$1I4621_DIB[6], _4I4657_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_766_5 (_4I4657_$1I4488_$1I4621_DIB[5], _4I4657_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_766_4 (_4I4657_$1I4488_$1I4621_DIB[4], _4I4657_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_766_3 (_4I4657_$1I4488_$1I4621_DIB[3], _4I4657_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_766_2 (_4I4657_$1I4488_$1I4621_DIB[2], _4I4657_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_766_1 (_4I4657_$1I4488_$1I4621_DIB[1], _4I4657_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_766_0 (_4I4657_$1I4488_$1I4621_DIB[0], _4I4657_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _4I4657_$1I4488_$1I4621_DIPA;
 reg [1:16] _4I4657_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_767_0 (_4I4657_$1I4488_$1I4621_DIPA[0], _4I4657_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _4I4657_$1I4488_$1I4621_DIPB;
 reg [1:16] _4I4657_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_768_1 (_4I4657_$1I4488_$1I4621_DIPB[1], _4I4657_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_768_0 (_4I4657_$1I4488_$1I4621_DIPB[0], _4I4657_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _4I4657_$1I4488_$1I4621_ENA;
 reg [1:16] _4I4657_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_769 (_4I4657_$1I4488_$1I4621_ENA, _4I4657_$1I4488_$1I4621_ENA__vlIN);

 wire  _4I4657_$1I4488_$1I4621_ENB;
 reg [1:16] _4I4657_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_770 (_4I4657_$1I4488_$1I4621_ENB, _4I4657_$1I4488_$1I4621_ENB__vlIN);

 wire  _4I4657_$1I4488_$1I4621_SSRA;
 reg [1:16] _4I4657_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_771 (_4I4657_$1I4488_$1I4621_SSRA, _4I4657_$1I4488_$1I4621_SSRA__vlIN);

 wire  _4I4657_$1I4488_$1I4621_SSRB;
 reg [1:16] _4I4657_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_772 (_4I4657_$1I4488_$1I4621_SSRB, _4I4657_$1I4488_$1I4621_SSRB__vlIN);

 wire  _4I4657_$1I4488_$1I4621_WEA;
 reg [1:16] _4I4657_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_773 (_4I4657_$1I4488_$1I4621_WEA, _4I4657_$1I4488_$1I4621_WEA__vlIN);

 wire  _4I4657_$1I4488_$1I4621_WEB;
 reg [1:16] _4I4657_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_774 (_4I4657_$1I4488_$1I4621_WEB, _4I4657_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _4I4657_$1I4488_$1I4621 ( _4I4657_$1I4488_$1I4621_DOA , _4I4657_$1I4488_$1I4621_DOB , _4I4657_$1I4488_$1I4621_DOPA , _4I4657_$1I4488_$1I4621_DOPB , _4I4657_$1I4488_$1I4621_ADDRA , _4I4657_$1I4488_$1I4621_ADDRB , _4I4657_$1I4488_$1I4621_CLKA , _4I4657_$1I4488_$1I4621_CLKB , _4I4657_$1I4488_$1I4621_DIA , _4I4657_$1I4488_$1I4621_DIB , _4I4657_$1I4488_$1I4621_DIPA , _4I4657_$1I4488_$1I4621_DIPB , _4I4657_$1I4488_$1I4621_ENA , _4I4657_$1I4488_$1I4621_ENB , _4I4657_$1I4488_$1I4621_SSRA , _4I4657_$1I4488_$1I4621_SSRB , _4I4657_$1I4488_$1I4621_WEA , _4I4657_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4657_$1I4488_$1I4620_DOA;

 wire [15:0] _4I4657_$1I4488_$1I4620_DOB;

 wire [0:0] _4I4657_$1I4488_$1I4620_DOPA;

 wire [1:0] _4I4657_$1I4488_$1I4620_DOPB;

 wire [10:0] _4I4657_$1I4488_$1I4620_ADDRA;
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_775_10 (_4I4657_$1I4488_$1I4620_ADDRA[10], _4I4657_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_775_9 (_4I4657_$1I4488_$1I4620_ADDRA[9], _4I4657_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_775_8 (_4I4657_$1I4488_$1I4620_ADDRA[8], _4I4657_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_775_7 (_4I4657_$1I4488_$1I4620_ADDRA[7], _4I4657_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_775_6 (_4I4657_$1I4488_$1I4620_ADDRA[6], _4I4657_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_775_5 (_4I4657_$1I4488_$1I4620_ADDRA[5], _4I4657_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_775_4 (_4I4657_$1I4488_$1I4620_ADDRA[4], _4I4657_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_775_3 (_4I4657_$1I4488_$1I4620_ADDRA[3], _4I4657_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_775_2 (_4I4657_$1I4488_$1I4620_ADDRA[2], _4I4657_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_775_1 (_4I4657_$1I4488_$1I4620_ADDRA[1], _4I4657_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_775_0 (_4I4657_$1I4488_$1I4620_ADDRA[0], _4I4657_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _4I4657_$1I4488_$1I4620_ADDRB;
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_776_9 (_4I4657_$1I4488_$1I4620_ADDRB[9], _4I4657_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_776_8 (_4I4657_$1I4488_$1I4620_ADDRB[8], _4I4657_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_776_7 (_4I4657_$1I4488_$1I4620_ADDRB[7], _4I4657_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_776_6 (_4I4657_$1I4488_$1I4620_ADDRB[6], _4I4657_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_776_5 (_4I4657_$1I4488_$1I4620_ADDRB[5], _4I4657_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_776_4 (_4I4657_$1I4488_$1I4620_ADDRB[4], _4I4657_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_776_3 (_4I4657_$1I4488_$1I4620_ADDRB[3], _4I4657_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_776_2 (_4I4657_$1I4488_$1I4620_ADDRB[2], _4I4657_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_776_1 (_4I4657_$1I4488_$1I4620_ADDRB[1], _4I4657_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_776_0 (_4I4657_$1I4488_$1I4620_ADDRB[0], _4I4657_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _4I4657_$1I4488_$1I4620_CLKA;
 reg [1:16] _4I4657_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_777 (_4I4657_$1I4488_$1I4620_CLKA, _4I4657_$1I4488_$1I4620_CLKA__vlIN);

 wire  _4I4657_$1I4488_$1I4620_CLKB;
 reg [1:16] _4I4657_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_778 (_4I4657_$1I4488_$1I4620_CLKB, _4I4657_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _4I4657_$1I4488_$1I4620_DIA;
 reg [1:16] _4I4657_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_779_7 (_4I4657_$1I4488_$1I4620_DIA[7], _4I4657_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_779_6 (_4I4657_$1I4488_$1I4620_DIA[6], _4I4657_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_779_5 (_4I4657_$1I4488_$1I4620_DIA[5], _4I4657_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_779_4 (_4I4657_$1I4488_$1I4620_DIA[4], _4I4657_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_779_3 (_4I4657_$1I4488_$1I4620_DIA[3], _4I4657_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_779_2 (_4I4657_$1I4488_$1I4620_DIA[2], _4I4657_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_779_1 (_4I4657_$1I4488_$1I4620_DIA[1], _4I4657_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_779_0 (_4I4657_$1I4488_$1I4620_DIA[0], _4I4657_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _4I4657_$1I4488_$1I4620_DIB;
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_780_15 (_4I4657_$1I4488_$1I4620_DIB[15], _4I4657_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_780_14 (_4I4657_$1I4488_$1I4620_DIB[14], _4I4657_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_780_13 (_4I4657_$1I4488_$1I4620_DIB[13], _4I4657_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_780_12 (_4I4657_$1I4488_$1I4620_DIB[12], _4I4657_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_780_11 (_4I4657_$1I4488_$1I4620_DIB[11], _4I4657_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_780_10 (_4I4657_$1I4488_$1I4620_DIB[10], _4I4657_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_780_9 (_4I4657_$1I4488_$1I4620_DIB[9], _4I4657_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_780_8 (_4I4657_$1I4488_$1I4620_DIB[8], _4I4657_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_780_7 (_4I4657_$1I4488_$1I4620_DIB[7], _4I4657_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_780_6 (_4I4657_$1I4488_$1I4620_DIB[6], _4I4657_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_780_5 (_4I4657_$1I4488_$1I4620_DIB[5], _4I4657_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_780_4 (_4I4657_$1I4488_$1I4620_DIB[4], _4I4657_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_780_3 (_4I4657_$1I4488_$1I4620_DIB[3], _4I4657_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_780_2 (_4I4657_$1I4488_$1I4620_DIB[2], _4I4657_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_780_1 (_4I4657_$1I4488_$1I4620_DIB[1], _4I4657_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_780_0 (_4I4657_$1I4488_$1I4620_DIB[0], _4I4657_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _4I4657_$1I4488_$1I4620_DIPA;
 reg [1:16] _4I4657_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_781_0 (_4I4657_$1I4488_$1I4620_DIPA[0], _4I4657_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _4I4657_$1I4488_$1I4620_DIPB;
 reg [1:16] _4I4657_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_782_1 (_4I4657_$1I4488_$1I4620_DIPB[1], _4I4657_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _4I4657_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_782_0 (_4I4657_$1I4488_$1I4620_DIPB[0], _4I4657_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _4I4657_$1I4488_$1I4620_ENA;
 reg [1:16] _4I4657_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_783 (_4I4657_$1I4488_$1I4620_ENA, _4I4657_$1I4488_$1I4620_ENA__vlIN);

 wire  _4I4657_$1I4488_$1I4620_ENB;
 reg [1:16] _4I4657_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_784 (_4I4657_$1I4488_$1I4620_ENB, _4I4657_$1I4488_$1I4620_ENB__vlIN);

 wire  _4I4657_$1I4488_$1I4620_SSRA;
 reg [1:16] _4I4657_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_785 (_4I4657_$1I4488_$1I4620_SSRA, _4I4657_$1I4488_$1I4620_SSRA__vlIN);

 wire  _4I4657_$1I4488_$1I4620_SSRB;
 reg [1:16] _4I4657_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_786 (_4I4657_$1I4488_$1I4620_SSRB, _4I4657_$1I4488_$1I4620_SSRB__vlIN);

 wire  _4I4657_$1I4488_$1I4620_WEA;
 reg [1:16] _4I4657_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_787 (_4I4657_$1I4488_$1I4620_WEA, _4I4657_$1I4488_$1I4620_WEA__vlIN);

 wire  _4I4657_$1I4488_$1I4620_WEB;
 reg [1:16] _4I4657_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_788 (_4I4657_$1I4488_$1I4620_WEB, _4I4657_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _4I4657_$1I4488_$1I4620 ( _4I4657_$1I4488_$1I4620_DOA , _4I4657_$1I4488_$1I4620_DOB , _4I4657_$1I4488_$1I4620_DOPA , _4I4657_$1I4488_$1I4620_DOPB , _4I4657_$1I4488_$1I4620_ADDRA , _4I4657_$1I4488_$1I4620_ADDRB , _4I4657_$1I4488_$1I4620_CLKA , _4I4657_$1I4488_$1I4620_CLKB , _4I4657_$1I4488_$1I4620_DIA , _4I4657_$1I4488_$1I4620_DIB , _4I4657_$1I4488_$1I4620_DIPA , _4I4657_$1I4488_$1I4620_DIPB , _4I4657_$1I4488_$1I4620_ENA , _4I4657_$1I4488_$1I4620_ENB , _4I4657_$1I4488_$1I4620_SSRA , _4I4657_$1I4488_$1I4620_SSRB , _4I4657_$1I4488_$1I4620_WEA , _4I4657_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4630_$1I4488_$1I4621_DOA;

 wire [15:0] _4I4630_$1I4488_$1I4621_DOB;

 wire [0:0] _4I4630_$1I4488_$1I4621_DOPA;

 wire [1:0] _4I4630_$1I4488_$1I4621_DOPB;

 wire [10:0] _4I4630_$1I4488_$1I4621_ADDRA;
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_789_10 (_4I4630_$1I4488_$1I4621_ADDRA[10], _4I4630_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_789_9 (_4I4630_$1I4488_$1I4621_ADDRA[9], _4I4630_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_789_8 (_4I4630_$1I4488_$1I4621_ADDRA[8], _4I4630_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_789_7 (_4I4630_$1I4488_$1I4621_ADDRA[7], _4I4630_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_789_6 (_4I4630_$1I4488_$1I4621_ADDRA[6], _4I4630_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_789_5 (_4I4630_$1I4488_$1I4621_ADDRA[5], _4I4630_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_789_4 (_4I4630_$1I4488_$1I4621_ADDRA[4], _4I4630_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_789_3 (_4I4630_$1I4488_$1I4621_ADDRA[3], _4I4630_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_789_2 (_4I4630_$1I4488_$1I4621_ADDRA[2], _4I4630_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_789_1 (_4I4630_$1I4488_$1I4621_ADDRA[1], _4I4630_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_789_0 (_4I4630_$1I4488_$1I4621_ADDRA[0], _4I4630_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _4I4630_$1I4488_$1I4621_ADDRB;
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_790_9 (_4I4630_$1I4488_$1I4621_ADDRB[9], _4I4630_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_790_8 (_4I4630_$1I4488_$1I4621_ADDRB[8], _4I4630_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_790_7 (_4I4630_$1I4488_$1I4621_ADDRB[7], _4I4630_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_790_6 (_4I4630_$1I4488_$1I4621_ADDRB[6], _4I4630_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_790_5 (_4I4630_$1I4488_$1I4621_ADDRB[5], _4I4630_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_790_4 (_4I4630_$1I4488_$1I4621_ADDRB[4], _4I4630_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_790_3 (_4I4630_$1I4488_$1I4621_ADDRB[3], _4I4630_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_790_2 (_4I4630_$1I4488_$1I4621_ADDRB[2], _4I4630_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_790_1 (_4I4630_$1I4488_$1I4621_ADDRB[1], _4I4630_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_790_0 (_4I4630_$1I4488_$1I4621_ADDRB[0], _4I4630_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _4I4630_$1I4488_$1I4621_CLKA;
 reg [1:16] _4I4630_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_791 (_4I4630_$1I4488_$1I4621_CLKA, _4I4630_$1I4488_$1I4621_CLKA__vlIN);

 wire  _4I4630_$1I4488_$1I4621_CLKB;
 reg [1:16] _4I4630_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_792 (_4I4630_$1I4488_$1I4621_CLKB, _4I4630_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _4I4630_$1I4488_$1I4621_DIA;
 reg [1:16] _4I4630_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_793_7 (_4I4630_$1I4488_$1I4621_DIA[7], _4I4630_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_793_6 (_4I4630_$1I4488_$1I4621_DIA[6], _4I4630_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_793_5 (_4I4630_$1I4488_$1I4621_DIA[5], _4I4630_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_793_4 (_4I4630_$1I4488_$1I4621_DIA[4], _4I4630_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_793_3 (_4I4630_$1I4488_$1I4621_DIA[3], _4I4630_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_793_2 (_4I4630_$1I4488_$1I4621_DIA[2], _4I4630_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_793_1 (_4I4630_$1I4488_$1I4621_DIA[1], _4I4630_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_793_0 (_4I4630_$1I4488_$1I4621_DIA[0], _4I4630_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _4I4630_$1I4488_$1I4621_DIB;
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_794_15 (_4I4630_$1I4488_$1I4621_DIB[15], _4I4630_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_794_14 (_4I4630_$1I4488_$1I4621_DIB[14], _4I4630_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_794_13 (_4I4630_$1I4488_$1I4621_DIB[13], _4I4630_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_794_12 (_4I4630_$1I4488_$1I4621_DIB[12], _4I4630_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_794_11 (_4I4630_$1I4488_$1I4621_DIB[11], _4I4630_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_794_10 (_4I4630_$1I4488_$1I4621_DIB[10], _4I4630_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_794_9 (_4I4630_$1I4488_$1I4621_DIB[9], _4I4630_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_794_8 (_4I4630_$1I4488_$1I4621_DIB[8], _4I4630_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_794_7 (_4I4630_$1I4488_$1I4621_DIB[7], _4I4630_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_794_6 (_4I4630_$1I4488_$1I4621_DIB[6], _4I4630_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_794_5 (_4I4630_$1I4488_$1I4621_DIB[5], _4I4630_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_794_4 (_4I4630_$1I4488_$1I4621_DIB[4], _4I4630_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_794_3 (_4I4630_$1I4488_$1I4621_DIB[3], _4I4630_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_794_2 (_4I4630_$1I4488_$1I4621_DIB[2], _4I4630_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_794_1 (_4I4630_$1I4488_$1I4621_DIB[1], _4I4630_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_794_0 (_4I4630_$1I4488_$1I4621_DIB[0], _4I4630_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _4I4630_$1I4488_$1I4621_DIPA;
 reg [1:16] _4I4630_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_795_0 (_4I4630_$1I4488_$1I4621_DIPA[0], _4I4630_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _4I4630_$1I4488_$1I4621_DIPB;
 reg [1:16] _4I4630_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_796_1 (_4I4630_$1I4488_$1I4621_DIPB[1], _4I4630_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_796_0 (_4I4630_$1I4488_$1I4621_DIPB[0], _4I4630_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _4I4630_$1I4488_$1I4621_ENA;
 reg [1:16] _4I4630_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_797 (_4I4630_$1I4488_$1I4621_ENA, _4I4630_$1I4488_$1I4621_ENA__vlIN);

 wire  _4I4630_$1I4488_$1I4621_ENB;
 reg [1:16] _4I4630_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_798 (_4I4630_$1I4488_$1I4621_ENB, _4I4630_$1I4488_$1I4621_ENB__vlIN);

 wire  _4I4630_$1I4488_$1I4621_SSRA;
 reg [1:16] _4I4630_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_799 (_4I4630_$1I4488_$1I4621_SSRA, _4I4630_$1I4488_$1I4621_SSRA__vlIN);

 wire  _4I4630_$1I4488_$1I4621_SSRB;
 reg [1:16] _4I4630_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_800 (_4I4630_$1I4488_$1I4621_SSRB, _4I4630_$1I4488_$1I4621_SSRB__vlIN);

 wire  _4I4630_$1I4488_$1I4621_WEA;
 reg [1:16] _4I4630_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_801 (_4I4630_$1I4488_$1I4621_WEA, _4I4630_$1I4488_$1I4621_WEA__vlIN);

 wire  _4I4630_$1I4488_$1I4621_WEB;
 reg [1:16] _4I4630_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_802 (_4I4630_$1I4488_$1I4621_WEB, _4I4630_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _4I4630_$1I4488_$1I4621 ( _4I4630_$1I4488_$1I4621_DOA , _4I4630_$1I4488_$1I4621_DOB , _4I4630_$1I4488_$1I4621_DOPA , _4I4630_$1I4488_$1I4621_DOPB , _4I4630_$1I4488_$1I4621_ADDRA , _4I4630_$1I4488_$1I4621_ADDRB , _4I4630_$1I4488_$1I4621_CLKA , _4I4630_$1I4488_$1I4621_CLKB , _4I4630_$1I4488_$1I4621_DIA , _4I4630_$1I4488_$1I4621_DIB , _4I4630_$1I4488_$1I4621_DIPA , _4I4630_$1I4488_$1I4621_DIPB , _4I4630_$1I4488_$1I4621_ENA , _4I4630_$1I4488_$1I4621_ENB , _4I4630_$1I4488_$1I4621_SSRA , _4I4630_$1I4488_$1I4621_SSRB , _4I4630_$1I4488_$1I4621_WEA , _4I4630_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4630_$1I4488_$1I4620_DOA;

 wire [15:0] _4I4630_$1I4488_$1I4620_DOB;

 wire [0:0] _4I4630_$1I4488_$1I4620_DOPA;

 wire [1:0] _4I4630_$1I4488_$1I4620_DOPB;

 wire [10:0] _4I4630_$1I4488_$1I4620_ADDRA;
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_803_10 (_4I4630_$1I4488_$1I4620_ADDRA[10], _4I4630_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_803_9 (_4I4630_$1I4488_$1I4620_ADDRA[9], _4I4630_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_803_8 (_4I4630_$1I4488_$1I4620_ADDRA[8], _4I4630_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_803_7 (_4I4630_$1I4488_$1I4620_ADDRA[7], _4I4630_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_803_6 (_4I4630_$1I4488_$1I4620_ADDRA[6], _4I4630_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_803_5 (_4I4630_$1I4488_$1I4620_ADDRA[5], _4I4630_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_803_4 (_4I4630_$1I4488_$1I4620_ADDRA[4], _4I4630_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_803_3 (_4I4630_$1I4488_$1I4620_ADDRA[3], _4I4630_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_803_2 (_4I4630_$1I4488_$1I4620_ADDRA[2], _4I4630_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_803_1 (_4I4630_$1I4488_$1I4620_ADDRA[1], _4I4630_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_803_0 (_4I4630_$1I4488_$1I4620_ADDRA[0], _4I4630_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _4I4630_$1I4488_$1I4620_ADDRB;
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_804_9 (_4I4630_$1I4488_$1I4620_ADDRB[9], _4I4630_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_804_8 (_4I4630_$1I4488_$1I4620_ADDRB[8], _4I4630_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_804_7 (_4I4630_$1I4488_$1I4620_ADDRB[7], _4I4630_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_804_6 (_4I4630_$1I4488_$1I4620_ADDRB[6], _4I4630_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_804_5 (_4I4630_$1I4488_$1I4620_ADDRB[5], _4I4630_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_804_4 (_4I4630_$1I4488_$1I4620_ADDRB[4], _4I4630_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_804_3 (_4I4630_$1I4488_$1I4620_ADDRB[3], _4I4630_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_804_2 (_4I4630_$1I4488_$1I4620_ADDRB[2], _4I4630_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_804_1 (_4I4630_$1I4488_$1I4620_ADDRB[1], _4I4630_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_804_0 (_4I4630_$1I4488_$1I4620_ADDRB[0], _4I4630_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _4I4630_$1I4488_$1I4620_CLKA;
 reg [1:16] _4I4630_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_805 (_4I4630_$1I4488_$1I4620_CLKA, _4I4630_$1I4488_$1I4620_CLKA__vlIN);

 wire  _4I4630_$1I4488_$1I4620_CLKB;
 reg [1:16] _4I4630_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_806 (_4I4630_$1I4488_$1I4620_CLKB, _4I4630_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _4I4630_$1I4488_$1I4620_DIA;
 reg [1:16] _4I4630_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_807_7 (_4I4630_$1I4488_$1I4620_DIA[7], _4I4630_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_807_6 (_4I4630_$1I4488_$1I4620_DIA[6], _4I4630_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_807_5 (_4I4630_$1I4488_$1I4620_DIA[5], _4I4630_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_807_4 (_4I4630_$1I4488_$1I4620_DIA[4], _4I4630_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_807_3 (_4I4630_$1I4488_$1I4620_DIA[3], _4I4630_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_807_2 (_4I4630_$1I4488_$1I4620_DIA[2], _4I4630_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_807_1 (_4I4630_$1I4488_$1I4620_DIA[1], _4I4630_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_807_0 (_4I4630_$1I4488_$1I4620_DIA[0], _4I4630_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _4I4630_$1I4488_$1I4620_DIB;
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_808_15 (_4I4630_$1I4488_$1I4620_DIB[15], _4I4630_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_808_14 (_4I4630_$1I4488_$1I4620_DIB[14], _4I4630_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_808_13 (_4I4630_$1I4488_$1I4620_DIB[13], _4I4630_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_808_12 (_4I4630_$1I4488_$1I4620_DIB[12], _4I4630_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_808_11 (_4I4630_$1I4488_$1I4620_DIB[11], _4I4630_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_808_10 (_4I4630_$1I4488_$1I4620_DIB[10], _4I4630_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_808_9 (_4I4630_$1I4488_$1I4620_DIB[9], _4I4630_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_808_8 (_4I4630_$1I4488_$1I4620_DIB[8], _4I4630_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_808_7 (_4I4630_$1I4488_$1I4620_DIB[7], _4I4630_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_808_6 (_4I4630_$1I4488_$1I4620_DIB[6], _4I4630_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_808_5 (_4I4630_$1I4488_$1I4620_DIB[5], _4I4630_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_808_4 (_4I4630_$1I4488_$1I4620_DIB[4], _4I4630_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_808_3 (_4I4630_$1I4488_$1I4620_DIB[3], _4I4630_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_808_2 (_4I4630_$1I4488_$1I4620_DIB[2], _4I4630_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_808_1 (_4I4630_$1I4488_$1I4620_DIB[1], _4I4630_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_808_0 (_4I4630_$1I4488_$1I4620_DIB[0], _4I4630_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _4I4630_$1I4488_$1I4620_DIPA;
 reg [1:16] _4I4630_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_809_0 (_4I4630_$1I4488_$1I4620_DIPA[0], _4I4630_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _4I4630_$1I4488_$1I4620_DIPB;
 reg [1:16] _4I4630_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_810_1 (_4I4630_$1I4488_$1I4620_DIPB[1], _4I4630_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _4I4630_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_810_0 (_4I4630_$1I4488_$1I4620_DIPB[0], _4I4630_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _4I4630_$1I4488_$1I4620_ENA;
 reg [1:16] _4I4630_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_811 (_4I4630_$1I4488_$1I4620_ENA, _4I4630_$1I4488_$1I4620_ENA__vlIN);

 wire  _4I4630_$1I4488_$1I4620_ENB;
 reg [1:16] _4I4630_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_812 (_4I4630_$1I4488_$1I4620_ENB, _4I4630_$1I4488_$1I4620_ENB__vlIN);

 wire  _4I4630_$1I4488_$1I4620_SSRA;
 reg [1:16] _4I4630_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_813 (_4I4630_$1I4488_$1I4620_SSRA, _4I4630_$1I4488_$1I4620_SSRA__vlIN);

 wire  _4I4630_$1I4488_$1I4620_SSRB;
 reg [1:16] _4I4630_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_814 (_4I4630_$1I4488_$1I4620_SSRB, _4I4630_$1I4488_$1I4620_SSRB__vlIN);

 wire  _4I4630_$1I4488_$1I4620_WEA;
 reg [1:16] _4I4630_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_815 (_4I4630_$1I4488_$1I4620_WEA, _4I4630_$1I4488_$1I4620_WEA__vlIN);

 wire  _4I4630_$1I4488_$1I4620_WEB;
 reg [1:16] _4I4630_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_816 (_4I4630_$1I4488_$1I4620_WEB, _4I4630_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _4I4630_$1I4488_$1I4620 ( _4I4630_$1I4488_$1I4620_DOA , _4I4630_$1I4488_$1I4620_DOB , _4I4630_$1I4488_$1I4620_DOPA , _4I4630_$1I4488_$1I4620_DOPB , _4I4630_$1I4488_$1I4620_ADDRA , _4I4630_$1I4488_$1I4620_ADDRB , _4I4630_$1I4488_$1I4620_CLKA , _4I4630_$1I4488_$1I4620_CLKB , _4I4630_$1I4488_$1I4620_DIA , _4I4630_$1I4488_$1I4620_DIB , _4I4630_$1I4488_$1I4620_DIPA , _4I4630_$1I4488_$1I4620_DIPB , _4I4630_$1I4488_$1I4620_ENA , _4I4630_$1I4488_$1I4620_ENB , _4I4630_$1I4488_$1I4620_SSRA , _4I4630_$1I4488_$1I4620_SSRB , _4I4630_$1I4488_$1I4620_WEA , _4I4630_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4611_$1I4488_$1I4621_DOA;

 wire [15:0] _4I4611_$1I4488_$1I4621_DOB;

 wire [0:0] _4I4611_$1I4488_$1I4621_DOPA;

 wire [1:0] _4I4611_$1I4488_$1I4621_DOPB;

 wire [10:0] _4I4611_$1I4488_$1I4621_ADDRA;
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_817_10 (_4I4611_$1I4488_$1I4621_ADDRA[10], _4I4611_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_817_9 (_4I4611_$1I4488_$1I4621_ADDRA[9], _4I4611_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_817_8 (_4I4611_$1I4488_$1I4621_ADDRA[8], _4I4611_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_817_7 (_4I4611_$1I4488_$1I4621_ADDRA[7], _4I4611_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_817_6 (_4I4611_$1I4488_$1I4621_ADDRA[6], _4I4611_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_817_5 (_4I4611_$1I4488_$1I4621_ADDRA[5], _4I4611_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_817_4 (_4I4611_$1I4488_$1I4621_ADDRA[4], _4I4611_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_817_3 (_4I4611_$1I4488_$1I4621_ADDRA[3], _4I4611_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_817_2 (_4I4611_$1I4488_$1I4621_ADDRA[2], _4I4611_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_817_1 (_4I4611_$1I4488_$1I4621_ADDRA[1], _4I4611_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_817_0 (_4I4611_$1I4488_$1I4621_ADDRA[0], _4I4611_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _4I4611_$1I4488_$1I4621_ADDRB;
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_818_9 (_4I4611_$1I4488_$1I4621_ADDRB[9], _4I4611_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_818_8 (_4I4611_$1I4488_$1I4621_ADDRB[8], _4I4611_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_818_7 (_4I4611_$1I4488_$1I4621_ADDRB[7], _4I4611_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_818_6 (_4I4611_$1I4488_$1I4621_ADDRB[6], _4I4611_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_818_5 (_4I4611_$1I4488_$1I4621_ADDRB[5], _4I4611_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_818_4 (_4I4611_$1I4488_$1I4621_ADDRB[4], _4I4611_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_818_3 (_4I4611_$1I4488_$1I4621_ADDRB[3], _4I4611_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_818_2 (_4I4611_$1I4488_$1I4621_ADDRB[2], _4I4611_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_818_1 (_4I4611_$1I4488_$1I4621_ADDRB[1], _4I4611_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_818_0 (_4I4611_$1I4488_$1I4621_ADDRB[0], _4I4611_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _4I4611_$1I4488_$1I4621_CLKA;
 reg [1:16] _4I4611_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_819 (_4I4611_$1I4488_$1I4621_CLKA, _4I4611_$1I4488_$1I4621_CLKA__vlIN);

 wire  _4I4611_$1I4488_$1I4621_CLKB;
 reg [1:16] _4I4611_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_820 (_4I4611_$1I4488_$1I4621_CLKB, _4I4611_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _4I4611_$1I4488_$1I4621_DIA;
 reg [1:16] _4I4611_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_821_7 (_4I4611_$1I4488_$1I4621_DIA[7], _4I4611_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_821_6 (_4I4611_$1I4488_$1I4621_DIA[6], _4I4611_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_821_5 (_4I4611_$1I4488_$1I4621_DIA[5], _4I4611_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_821_4 (_4I4611_$1I4488_$1I4621_DIA[4], _4I4611_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_821_3 (_4I4611_$1I4488_$1I4621_DIA[3], _4I4611_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_821_2 (_4I4611_$1I4488_$1I4621_DIA[2], _4I4611_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_821_1 (_4I4611_$1I4488_$1I4621_DIA[1], _4I4611_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_821_0 (_4I4611_$1I4488_$1I4621_DIA[0], _4I4611_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _4I4611_$1I4488_$1I4621_DIB;
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_822_15 (_4I4611_$1I4488_$1I4621_DIB[15], _4I4611_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_822_14 (_4I4611_$1I4488_$1I4621_DIB[14], _4I4611_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_822_13 (_4I4611_$1I4488_$1I4621_DIB[13], _4I4611_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_822_12 (_4I4611_$1I4488_$1I4621_DIB[12], _4I4611_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_822_11 (_4I4611_$1I4488_$1I4621_DIB[11], _4I4611_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_822_10 (_4I4611_$1I4488_$1I4621_DIB[10], _4I4611_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_822_9 (_4I4611_$1I4488_$1I4621_DIB[9], _4I4611_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_822_8 (_4I4611_$1I4488_$1I4621_DIB[8], _4I4611_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_822_7 (_4I4611_$1I4488_$1I4621_DIB[7], _4I4611_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_822_6 (_4I4611_$1I4488_$1I4621_DIB[6], _4I4611_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_822_5 (_4I4611_$1I4488_$1I4621_DIB[5], _4I4611_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_822_4 (_4I4611_$1I4488_$1I4621_DIB[4], _4I4611_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_822_3 (_4I4611_$1I4488_$1I4621_DIB[3], _4I4611_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_822_2 (_4I4611_$1I4488_$1I4621_DIB[2], _4I4611_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_822_1 (_4I4611_$1I4488_$1I4621_DIB[1], _4I4611_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_822_0 (_4I4611_$1I4488_$1I4621_DIB[0], _4I4611_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _4I4611_$1I4488_$1I4621_DIPA;
 reg [1:16] _4I4611_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_823_0 (_4I4611_$1I4488_$1I4621_DIPA[0], _4I4611_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _4I4611_$1I4488_$1I4621_DIPB;
 reg [1:16] _4I4611_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_824_1 (_4I4611_$1I4488_$1I4621_DIPB[1], _4I4611_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_824_0 (_4I4611_$1I4488_$1I4621_DIPB[0], _4I4611_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _4I4611_$1I4488_$1I4621_ENA;
 reg [1:16] _4I4611_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_825 (_4I4611_$1I4488_$1I4621_ENA, _4I4611_$1I4488_$1I4621_ENA__vlIN);

 wire  _4I4611_$1I4488_$1I4621_ENB;
 reg [1:16] _4I4611_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_826 (_4I4611_$1I4488_$1I4621_ENB, _4I4611_$1I4488_$1I4621_ENB__vlIN);

 wire  _4I4611_$1I4488_$1I4621_SSRA;
 reg [1:16] _4I4611_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_827 (_4I4611_$1I4488_$1I4621_SSRA, _4I4611_$1I4488_$1I4621_SSRA__vlIN);

 wire  _4I4611_$1I4488_$1I4621_SSRB;
 reg [1:16] _4I4611_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_828 (_4I4611_$1I4488_$1I4621_SSRB, _4I4611_$1I4488_$1I4621_SSRB__vlIN);

 wire  _4I4611_$1I4488_$1I4621_WEA;
 reg [1:16] _4I4611_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_829 (_4I4611_$1I4488_$1I4621_WEA, _4I4611_$1I4488_$1I4621_WEA__vlIN);

 wire  _4I4611_$1I4488_$1I4621_WEB;
 reg [1:16] _4I4611_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_830 (_4I4611_$1I4488_$1I4621_WEB, _4I4611_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _4I4611_$1I4488_$1I4621 ( _4I4611_$1I4488_$1I4621_DOA , _4I4611_$1I4488_$1I4621_DOB , _4I4611_$1I4488_$1I4621_DOPA , _4I4611_$1I4488_$1I4621_DOPB , _4I4611_$1I4488_$1I4621_ADDRA , _4I4611_$1I4488_$1I4621_ADDRB , _4I4611_$1I4488_$1I4621_CLKA , _4I4611_$1I4488_$1I4621_CLKB , _4I4611_$1I4488_$1I4621_DIA , _4I4611_$1I4488_$1I4621_DIB , _4I4611_$1I4488_$1I4621_DIPA , _4I4611_$1I4488_$1I4621_DIPB , _4I4611_$1I4488_$1I4621_ENA , _4I4611_$1I4488_$1I4621_ENB , _4I4611_$1I4488_$1I4621_SSRA , _4I4611_$1I4488_$1I4621_SSRB , _4I4611_$1I4488_$1I4621_WEA , _4I4611_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4611_$1I4488_$1I4620_DOA;

 wire [15:0] _4I4611_$1I4488_$1I4620_DOB;

 wire [0:0] _4I4611_$1I4488_$1I4620_DOPA;

 wire [1:0] _4I4611_$1I4488_$1I4620_DOPB;

 wire [10:0] _4I4611_$1I4488_$1I4620_ADDRA;
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_831_10 (_4I4611_$1I4488_$1I4620_ADDRA[10], _4I4611_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_831_9 (_4I4611_$1I4488_$1I4620_ADDRA[9], _4I4611_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_831_8 (_4I4611_$1I4488_$1I4620_ADDRA[8], _4I4611_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_831_7 (_4I4611_$1I4488_$1I4620_ADDRA[7], _4I4611_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_831_6 (_4I4611_$1I4488_$1I4620_ADDRA[6], _4I4611_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_831_5 (_4I4611_$1I4488_$1I4620_ADDRA[5], _4I4611_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_831_4 (_4I4611_$1I4488_$1I4620_ADDRA[4], _4I4611_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_831_3 (_4I4611_$1I4488_$1I4620_ADDRA[3], _4I4611_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_831_2 (_4I4611_$1I4488_$1I4620_ADDRA[2], _4I4611_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_831_1 (_4I4611_$1I4488_$1I4620_ADDRA[1], _4I4611_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_831_0 (_4I4611_$1I4488_$1I4620_ADDRA[0], _4I4611_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _4I4611_$1I4488_$1I4620_ADDRB;
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_832_9 (_4I4611_$1I4488_$1I4620_ADDRB[9], _4I4611_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_832_8 (_4I4611_$1I4488_$1I4620_ADDRB[8], _4I4611_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_832_7 (_4I4611_$1I4488_$1I4620_ADDRB[7], _4I4611_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_832_6 (_4I4611_$1I4488_$1I4620_ADDRB[6], _4I4611_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_832_5 (_4I4611_$1I4488_$1I4620_ADDRB[5], _4I4611_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_832_4 (_4I4611_$1I4488_$1I4620_ADDRB[4], _4I4611_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_832_3 (_4I4611_$1I4488_$1I4620_ADDRB[3], _4I4611_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_832_2 (_4I4611_$1I4488_$1I4620_ADDRB[2], _4I4611_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_832_1 (_4I4611_$1I4488_$1I4620_ADDRB[1], _4I4611_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_832_0 (_4I4611_$1I4488_$1I4620_ADDRB[0], _4I4611_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _4I4611_$1I4488_$1I4620_CLKA;
 reg [1:16] _4I4611_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_833 (_4I4611_$1I4488_$1I4620_CLKA, _4I4611_$1I4488_$1I4620_CLKA__vlIN);

 wire  _4I4611_$1I4488_$1I4620_CLKB;
 reg [1:16] _4I4611_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_834 (_4I4611_$1I4488_$1I4620_CLKB, _4I4611_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _4I4611_$1I4488_$1I4620_DIA;
 reg [1:16] _4I4611_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_835_7 (_4I4611_$1I4488_$1I4620_DIA[7], _4I4611_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_835_6 (_4I4611_$1I4488_$1I4620_DIA[6], _4I4611_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_835_5 (_4I4611_$1I4488_$1I4620_DIA[5], _4I4611_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_835_4 (_4I4611_$1I4488_$1I4620_DIA[4], _4I4611_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_835_3 (_4I4611_$1I4488_$1I4620_DIA[3], _4I4611_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_835_2 (_4I4611_$1I4488_$1I4620_DIA[2], _4I4611_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_835_1 (_4I4611_$1I4488_$1I4620_DIA[1], _4I4611_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_835_0 (_4I4611_$1I4488_$1I4620_DIA[0], _4I4611_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _4I4611_$1I4488_$1I4620_DIB;
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_836_15 (_4I4611_$1I4488_$1I4620_DIB[15], _4I4611_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_836_14 (_4I4611_$1I4488_$1I4620_DIB[14], _4I4611_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_836_13 (_4I4611_$1I4488_$1I4620_DIB[13], _4I4611_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_836_12 (_4I4611_$1I4488_$1I4620_DIB[12], _4I4611_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_836_11 (_4I4611_$1I4488_$1I4620_DIB[11], _4I4611_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_836_10 (_4I4611_$1I4488_$1I4620_DIB[10], _4I4611_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_836_9 (_4I4611_$1I4488_$1I4620_DIB[9], _4I4611_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_836_8 (_4I4611_$1I4488_$1I4620_DIB[8], _4I4611_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_836_7 (_4I4611_$1I4488_$1I4620_DIB[7], _4I4611_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_836_6 (_4I4611_$1I4488_$1I4620_DIB[6], _4I4611_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_836_5 (_4I4611_$1I4488_$1I4620_DIB[5], _4I4611_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_836_4 (_4I4611_$1I4488_$1I4620_DIB[4], _4I4611_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_836_3 (_4I4611_$1I4488_$1I4620_DIB[3], _4I4611_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_836_2 (_4I4611_$1I4488_$1I4620_DIB[2], _4I4611_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_836_1 (_4I4611_$1I4488_$1I4620_DIB[1], _4I4611_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_836_0 (_4I4611_$1I4488_$1I4620_DIB[0], _4I4611_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _4I4611_$1I4488_$1I4620_DIPA;
 reg [1:16] _4I4611_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_837_0 (_4I4611_$1I4488_$1I4620_DIPA[0], _4I4611_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _4I4611_$1I4488_$1I4620_DIPB;
 reg [1:16] _4I4611_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_838_1 (_4I4611_$1I4488_$1I4620_DIPB[1], _4I4611_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _4I4611_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_838_0 (_4I4611_$1I4488_$1I4620_DIPB[0], _4I4611_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _4I4611_$1I4488_$1I4620_ENA;
 reg [1:16] _4I4611_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_839 (_4I4611_$1I4488_$1I4620_ENA, _4I4611_$1I4488_$1I4620_ENA__vlIN);

 wire  _4I4611_$1I4488_$1I4620_ENB;
 reg [1:16] _4I4611_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_840 (_4I4611_$1I4488_$1I4620_ENB, _4I4611_$1I4488_$1I4620_ENB__vlIN);

 wire  _4I4611_$1I4488_$1I4620_SSRA;
 reg [1:16] _4I4611_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_841 (_4I4611_$1I4488_$1I4620_SSRA, _4I4611_$1I4488_$1I4620_SSRA__vlIN);

 wire  _4I4611_$1I4488_$1I4620_SSRB;
 reg [1:16] _4I4611_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_842 (_4I4611_$1I4488_$1I4620_SSRB, _4I4611_$1I4488_$1I4620_SSRB__vlIN);

 wire  _4I4611_$1I4488_$1I4620_WEA;
 reg [1:16] _4I4611_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_843 (_4I4611_$1I4488_$1I4620_WEA, _4I4611_$1I4488_$1I4620_WEA__vlIN);

 wire  _4I4611_$1I4488_$1I4620_WEB;
 reg [1:16] _4I4611_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_844 (_4I4611_$1I4488_$1I4620_WEB, _4I4611_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _4I4611_$1I4488_$1I4620 ( _4I4611_$1I4488_$1I4620_DOA , _4I4611_$1I4488_$1I4620_DOB , _4I4611_$1I4488_$1I4620_DOPA , _4I4611_$1I4488_$1I4620_DOPB , _4I4611_$1I4488_$1I4620_ADDRA , _4I4611_$1I4488_$1I4620_ADDRB , _4I4611_$1I4488_$1I4620_CLKA , _4I4611_$1I4488_$1I4620_CLKB , _4I4611_$1I4488_$1I4620_DIA , _4I4611_$1I4488_$1I4620_DIB , _4I4611_$1I4488_$1I4620_DIPA , _4I4611_$1I4488_$1I4620_DIPB , _4I4611_$1I4488_$1I4620_ENA , _4I4611_$1I4488_$1I4620_ENB , _4I4611_$1I4488_$1I4620_SSRA , _4I4611_$1I4488_$1I4620_SSRB , _4I4611_$1I4488_$1I4620_WEA , _4I4611_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4560_$1I4488_$1I4621_DOA;

 wire [15:0] _4I4560_$1I4488_$1I4621_DOB;

 wire [0:0] _4I4560_$1I4488_$1I4621_DOPA;

 wire [1:0] _4I4560_$1I4488_$1I4621_DOPB;

 wire [10:0] _4I4560_$1I4488_$1I4621_ADDRA;
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_845_10 (_4I4560_$1I4488_$1I4621_ADDRA[10], _4I4560_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_845_9 (_4I4560_$1I4488_$1I4621_ADDRA[9], _4I4560_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_845_8 (_4I4560_$1I4488_$1I4621_ADDRA[8], _4I4560_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_845_7 (_4I4560_$1I4488_$1I4621_ADDRA[7], _4I4560_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_845_6 (_4I4560_$1I4488_$1I4621_ADDRA[6], _4I4560_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_845_5 (_4I4560_$1I4488_$1I4621_ADDRA[5], _4I4560_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_845_4 (_4I4560_$1I4488_$1I4621_ADDRA[4], _4I4560_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_845_3 (_4I4560_$1I4488_$1I4621_ADDRA[3], _4I4560_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_845_2 (_4I4560_$1I4488_$1I4621_ADDRA[2], _4I4560_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_845_1 (_4I4560_$1I4488_$1I4621_ADDRA[1], _4I4560_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_845_0 (_4I4560_$1I4488_$1I4621_ADDRA[0], _4I4560_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _4I4560_$1I4488_$1I4621_ADDRB;
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_846_9 (_4I4560_$1I4488_$1I4621_ADDRB[9], _4I4560_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_846_8 (_4I4560_$1I4488_$1I4621_ADDRB[8], _4I4560_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_846_7 (_4I4560_$1I4488_$1I4621_ADDRB[7], _4I4560_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_846_6 (_4I4560_$1I4488_$1I4621_ADDRB[6], _4I4560_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_846_5 (_4I4560_$1I4488_$1I4621_ADDRB[5], _4I4560_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_846_4 (_4I4560_$1I4488_$1I4621_ADDRB[4], _4I4560_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_846_3 (_4I4560_$1I4488_$1I4621_ADDRB[3], _4I4560_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_846_2 (_4I4560_$1I4488_$1I4621_ADDRB[2], _4I4560_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_846_1 (_4I4560_$1I4488_$1I4621_ADDRB[1], _4I4560_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_846_0 (_4I4560_$1I4488_$1I4621_ADDRB[0], _4I4560_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _4I4560_$1I4488_$1I4621_CLKA;
 reg [1:16] _4I4560_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_847 (_4I4560_$1I4488_$1I4621_CLKA, _4I4560_$1I4488_$1I4621_CLKA__vlIN);

 wire  _4I4560_$1I4488_$1I4621_CLKB;
 reg [1:16] _4I4560_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_848 (_4I4560_$1I4488_$1I4621_CLKB, _4I4560_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _4I4560_$1I4488_$1I4621_DIA;
 reg [1:16] _4I4560_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_849_7 (_4I4560_$1I4488_$1I4621_DIA[7], _4I4560_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_849_6 (_4I4560_$1I4488_$1I4621_DIA[6], _4I4560_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_849_5 (_4I4560_$1I4488_$1I4621_DIA[5], _4I4560_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_849_4 (_4I4560_$1I4488_$1I4621_DIA[4], _4I4560_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_849_3 (_4I4560_$1I4488_$1I4621_DIA[3], _4I4560_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_849_2 (_4I4560_$1I4488_$1I4621_DIA[2], _4I4560_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_849_1 (_4I4560_$1I4488_$1I4621_DIA[1], _4I4560_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_849_0 (_4I4560_$1I4488_$1I4621_DIA[0], _4I4560_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _4I4560_$1I4488_$1I4621_DIB;
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_850_15 (_4I4560_$1I4488_$1I4621_DIB[15], _4I4560_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_850_14 (_4I4560_$1I4488_$1I4621_DIB[14], _4I4560_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_850_13 (_4I4560_$1I4488_$1I4621_DIB[13], _4I4560_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_850_12 (_4I4560_$1I4488_$1I4621_DIB[12], _4I4560_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_850_11 (_4I4560_$1I4488_$1I4621_DIB[11], _4I4560_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_850_10 (_4I4560_$1I4488_$1I4621_DIB[10], _4I4560_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_850_9 (_4I4560_$1I4488_$1I4621_DIB[9], _4I4560_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_850_8 (_4I4560_$1I4488_$1I4621_DIB[8], _4I4560_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_850_7 (_4I4560_$1I4488_$1I4621_DIB[7], _4I4560_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_850_6 (_4I4560_$1I4488_$1I4621_DIB[6], _4I4560_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_850_5 (_4I4560_$1I4488_$1I4621_DIB[5], _4I4560_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_850_4 (_4I4560_$1I4488_$1I4621_DIB[4], _4I4560_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_850_3 (_4I4560_$1I4488_$1I4621_DIB[3], _4I4560_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_850_2 (_4I4560_$1I4488_$1I4621_DIB[2], _4I4560_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_850_1 (_4I4560_$1I4488_$1I4621_DIB[1], _4I4560_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_850_0 (_4I4560_$1I4488_$1I4621_DIB[0], _4I4560_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _4I4560_$1I4488_$1I4621_DIPA;
 reg [1:16] _4I4560_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_851_0 (_4I4560_$1I4488_$1I4621_DIPA[0], _4I4560_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _4I4560_$1I4488_$1I4621_DIPB;
 reg [1:16] _4I4560_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_852_1 (_4I4560_$1I4488_$1I4621_DIPB[1], _4I4560_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_852_0 (_4I4560_$1I4488_$1I4621_DIPB[0], _4I4560_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _4I4560_$1I4488_$1I4621_ENA;
 reg [1:16] _4I4560_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_853 (_4I4560_$1I4488_$1I4621_ENA, _4I4560_$1I4488_$1I4621_ENA__vlIN);

 wire  _4I4560_$1I4488_$1I4621_ENB;
 reg [1:16] _4I4560_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_854 (_4I4560_$1I4488_$1I4621_ENB, _4I4560_$1I4488_$1I4621_ENB__vlIN);

 wire  _4I4560_$1I4488_$1I4621_SSRA;
 reg [1:16] _4I4560_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_855 (_4I4560_$1I4488_$1I4621_SSRA, _4I4560_$1I4488_$1I4621_SSRA__vlIN);

 wire  _4I4560_$1I4488_$1I4621_SSRB;
 reg [1:16] _4I4560_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_856 (_4I4560_$1I4488_$1I4621_SSRB, _4I4560_$1I4488_$1I4621_SSRB__vlIN);

 wire  _4I4560_$1I4488_$1I4621_WEA;
 reg [1:16] _4I4560_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_857 (_4I4560_$1I4488_$1I4621_WEA, _4I4560_$1I4488_$1I4621_WEA__vlIN);

 wire  _4I4560_$1I4488_$1I4621_WEB;
 reg [1:16] _4I4560_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_858 (_4I4560_$1I4488_$1I4621_WEB, _4I4560_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _4I4560_$1I4488_$1I4621 ( _4I4560_$1I4488_$1I4621_DOA , _4I4560_$1I4488_$1I4621_DOB , _4I4560_$1I4488_$1I4621_DOPA , _4I4560_$1I4488_$1I4621_DOPB , _4I4560_$1I4488_$1I4621_ADDRA , _4I4560_$1I4488_$1I4621_ADDRB , _4I4560_$1I4488_$1I4621_CLKA , _4I4560_$1I4488_$1I4621_CLKB , _4I4560_$1I4488_$1I4621_DIA , _4I4560_$1I4488_$1I4621_DIB , _4I4560_$1I4488_$1I4621_DIPA , _4I4560_$1I4488_$1I4621_DIPB , _4I4560_$1I4488_$1I4621_ENA , _4I4560_$1I4488_$1I4621_ENB , _4I4560_$1I4488_$1I4621_SSRA , _4I4560_$1I4488_$1I4621_SSRB , _4I4560_$1I4488_$1I4621_WEA , _4I4560_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4560_$1I4488_$1I4620_DOA;

 wire [15:0] _4I4560_$1I4488_$1I4620_DOB;

 wire [0:0] _4I4560_$1I4488_$1I4620_DOPA;

 wire [1:0] _4I4560_$1I4488_$1I4620_DOPB;

 wire [10:0] _4I4560_$1I4488_$1I4620_ADDRA;
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_859_10 (_4I4560_$1I4488_$1I4620_ADDRA[10], _4I4560_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_859_9 (_4I4560_$1I4488_$1I4620_ADDRA[9], _4I4560_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_859_8 (_4I4560_$1I4488_$1I4620_ADDRA[8], _4I4560_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_859_7 (_4I4560_$1I4488_$1I4620_ADDRA[7], _4I4560_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_859_6 (_4I4560_$1I4488_$1I4620_ADDRA[6], _4I4560_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_859_5 (_4I4560_$1I4488_$1I4620_ADDRA[5], _4I4560_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_859_4 (_4I4560_$1I4488_$1I4620_ADDRA[4], _4I4560_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_859_3 (_4I4560_$1I4488_$1I4620_ADDRA[3], _4I4560_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_859_2 (_4I4560_$1I4488_$1I4620_ADDRA[2], _4I4560_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_859_1 (_4I4560_$1I4488_$1I4620_ADDRA[1], _4I4560_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_859_0 (_4I4560_$1I4488_$1I4620_ADDRA[0], _4I4560_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _4I4560_$1I4488_$1I4620_ADDRB;
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_860_9 (_4I4560_$1I4488_$1I4620_ADDRB[9], _4I4560_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_860_8 (_4I4560_$1I4488_$1I4620_ADDRB[8], _4I4560_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_860_7 (_4I4560_$1I4488_$1I4620_ADDRB[7], _4I4560_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_860_6 (_4I4560_$1I4488_$1I4620_ADDRB[6], _4I4560_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_860_5 (_4I4560_$1I4488_$1I4620_ADDRB[5], _4I4560_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_860_4 (_4I4560_$1I4488_$1I4620_ADDRB[4], _4I4560_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_860_3 (_4I4560_$1I4488_$1I4620_ADDRB[3], _4I4560_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_860_2 (_4I4560_$1I4488_$1I4620_ADDRB[2], _4I4560_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_860_1 (_4I4560_$1I4488_$1I4620_ADDRB[1], _4I4560_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_860_0 (_4I4560_$1I4488_$1I4620_ADDRB[0], _4I4560_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _4I4560_$1I4488_$1I4620_CLKA;
 reg [1:16] _4I4560_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_861 (_4I4560_$1I4488_$1I4620_CLKA, _4I4560_$1I4488_$1I4620_CLKA__vlIN);

 wire  _4I4560_$1I4488_$1I4620_CLKB;
 reg [1:16] _4I4560_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_862 (_4I4560_$1I4488_$1I4620_CLKB, _4I4560_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _4I4560_$1I4488_$1I4620_DIA;
 reg [1:16] _4I4560_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_863_7 (_4I4560_$1I4488_$1I4620_DIA[7], _4I4560_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_863_6 (_4I4560_$1I4488_$1I4620_DIA[6], _4I4560_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_863_5 (_4I4560_$1I4488_$1I4620_DIA[5], _4I4560_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_863_4 (_4I4560_$1I4488_$1I4620_DIA[4], _4I4560_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_863_3 (_4I4560_$1I4488_$1I4620_DIA[3], _4I4560_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_863_2 (_4I4560_$1I4488_$1I4620_DIA[2], _4I4560_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_863_1 (_4I4560_$1I4488_$1I4620_DIA[1], _4I4560_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_863_0 (_4I4560_$1I4488_$1I4620_DIA[0], _4I4560_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _4I4560_$1I4488_$1I4620_DIB;
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_864_15 (_4I4560_$1I4488_$1I4620_DIB[15], _4I4560_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_864_14 (_4I4560_$1I4488_$1I4620_DIB[14], _4I4560_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_864_13 (_4I4560_$1I4488_$1I4620_DIB[13], _4I4560_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_864_12 (_4I4560_$1I4488_$1I4620_DIB[12], _4I4560_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_864_11 (_4I4560_$1I4488_$1I4620_DIB[11], _4I4560_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_864_10 (_4I4560_$1I4488_$1I4620_DIB[10], _4I4560_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_864_9 (_4I4560_$1I4488_$1I4620_DIB[9], _4I4560_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_864_8 (_4I4560_$1I4488_$1I4620_DIB[8], _4I4560_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_864_7 (_4I4560_$1I4488_$1I4620_DIB[7], _4I4560_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_864_6 (_4I4560_$1I4488_$1I4620_DIB[6], _4I4560_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_864_5 (_4I4560_$1I4488_$1I4620_DIB[5], _4I4560_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_864_4 (_4I4560_$1I4488_$1I4620_DIB[4], _4I4560_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_864_3 (_4I4560_$1I4488_$1I4620_DIB[3], _4I4560_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_864_2 (_4I4560_$1I4488_$1I4620_DIB[2], _4I4560_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_864_1 (_4I4560_$1I4488_$1I4620_DIB[1], _4I4560_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_864_0 (_4I4560_$1I4488_$1I4620_DIB[0], _4I4560_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _4I4560_$1I4488_$1I4620_DIPA;
 reg [1:16] _4I4560_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_865_0 (_4I4560_$1I4488_$1I4620_DIPA[0], _4I4560_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _4I4560_$1I4488_$1I4620_DIPB;
 reg [1:16] _4I4560_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_866_1 (_4I4560_$1I4488_$1I4620_DIPB[1], _4I4560_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _4I4560_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_866_0 (_4I4560_$1I4488_$1I4620_DIPB[0], _4I4560_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _4I4560_$1I4488_$1I4620_ENA;
 reg [1:16] _4I4560_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_867 (_4I4560_$1I4488_$1I4620_ENA, _4I4560_$1I4488_$1I4620_ENA__vlIN);

 wire  _4I4560_$1I4488_$1I4620_ENB;
 reg [1:16] _4I4560_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_868 (_4I4560_$1I4488_$1I4620_ENB, _4I4560_$1I4488_$1I4620_ENB__vlIN);

 wire  _4I4560_$1I4488_$1I4620_SSRA;
 reg [1:16] _4I4560_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_869 (_4I4560_$1I4488_$1I4620_SSRA, _4I4560_$1I4488_$1I4620_SSRA__vlIN);

 wire  _4I4560_$1I4488_$1I4620_SSRB;
 reg [1:16] _4I4560_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_870 (_4I4560_$1I4488_$1I4620_SSRB, _4I4560_$1I4488_$1I4620_SSRB__vlIN);

 wire  _4I4560_$1I4488_$1I4620_WEA;
 reg [1:16] _4I4560_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_871 (_4I4560_$1I4488_$1I4620_WEA, _4I4560_$1I4488_$1I4620_WEA__vlIN);

 wire  _4I4560_$1I4488_$1I4620_WEB;
 reg [1:16] _4I4560_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_872 (_4I4560_$1I4488_$1I4620_WEB, _4I4560_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _4I4560_$1I4488_$1I4620 ( _4I4560_$1I4488_$1I4620_DOA , _4I4560_$1I4488_$1I4620_DOB , _4I4560_$1I4488_$1I4620_DOPA , _4I4560_$1I4488_$1I4620_DOPB , _4I4560_$1I4488_$1I4620_ADDRA , _4I4560_$1I4488_$1I4620_ADDRB , _4I4560_$1I4488_$1I4620_CLKA , _4I4560_$1I4488_$1I4620_CLKB , _4I4560_$1I4488_$1I4620_DIA , _4I4560_$1I4488_$1I4620_DIB , _4I4560_$1I4488_$1I4620_DIPA , _4I4560_$1I4488_$1I4620_DIPB , _4I4560_$1I4488_$1I4620_ENA , _4I4560_$1I4488_$1I4620_ENB , _4I4560_$1I4488_$1I4620_SSRA , _4I4560_$1I4488_$1I4620_SSRB , _4I4560_$1I4488_$1I4620_WEA , _4I4560_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4526_$1I4488_$1I4621_DOA;

 wire [15:0] _4I4526_$1I4488_$1I4621_DOB;

 wire [0:0] _4I4526_$1I4488_$1I4621_DOPA;

 wire [1:0] _4I4526_$1I4488_$1I4621_DOPB;

 wire [10:0] _4I4526_$1I4488_$1I4621_ADDRA;
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_873_10 (_4I4526_$1I4488_$1I4621_ADDRA[10], _4I4526_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_873_9 (_4I4526_$1I4488_$1I4621_ADDRA[9], _4I4526_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_873_8 (_4I4526_$1I4488_$1I4621_ADDRA[8], _4I4526_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_873_7 (_4I4526_$1I4488_$1I4621_ADDRA[7], _4I4526_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_873_6 (_4I4526_$1I4488_$1I4621_ADDRA[6], _4I4526_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_873_5 (_4I4526_$1I4488_$1I4621_ADDRA[5], _4I4526_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_873_4 (_4I4526_$1I4488_$1I4621_ADDRA[4], _4I4526_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_873_3 (_4I4526_$1I4488_$1I4621_ADDRA[3], _4I4526_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_873_2 (_4I4526_$1I4488_$1I4621_ADDRA[2], _4I4526_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_873_1 (_4I4526_$1I4488_$1I4621_ADDRA[1], _4I4526_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_873_0 (_4I4526_$1I4488_$1I4621_ADDRA[0], _4I4526_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _4I4526_$1I4488_$1I4621_ADDRB;
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_874_9 (_4I4526_$1I4488_$1I4621_ADDRB[9], _4I4526_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_874_8 (_4I4526_$1I4488_$1I4621_ADDRB[8], _4I4526_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_874_7 (_4I4526_$1I4488_$1I4621_ADDRB[7], _4I4526_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_874_6 (_4I4526_$1I4488_$1I4621_ADDRB[6], _4I4526_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_874_5 (_4I4526_$1I4488_$1I4621_ADDRB[5], _4I4526_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_874_4 (_4I4526_$1I4488_$1I4621_ADDRB[4], _4I4526_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_874_3 (_4I4526_$1I4488_$1I4621_ADDRB[3], _4I4526_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_874_2 (_4I4526_$1I4488_$1I4621_ADDRB[2], _4I4526_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_874_1 (_4I4526_$1I4488_$1I4621_ADDRB[1], _4I4526_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_874_0 (_4I4526_$1I4488_$1I4621_ADDRB[0], _4I4526_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _4I4526_$1I4488_$1I4621_CLKA;
 reg [1:16] _4I4526_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_875 (_4I4526_$1I4488_$1I4621_CLKA, _4I4526_$1I4488_$1I4621_CLKA__vlIN);

 wire  _4I4526_$1I4488_$1I4621_CLKB;
 reg [1:16] _4I4526_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_876 (_4I4526_$1I4488_$1I4621_CLKB, _4I4526_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _4I4526_$1I4488_$1I4621_DIA;
 reg [1:16] _4I4526_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_877_7 (_4I4526_$1I4488_$1I4621_DIA[7], _4I4526_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_877_6 (_4I4526_$1I4488_$1I4621_DIA[6], _4I4526_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_877_5 (_4I4526_$1I4488_$1I4621_DIA[5], _4I4526_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_877_4 (_4I4526_$1I4488_$1I4621_DIA[4], _4I4526_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_877_3 (_4I4526_$1I4488_$1I4621_DIA[3], _4I4526_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_877_2 (_4I4526_$1I4488_$1I4621_DIA[2], _4I4526_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_877_1 (_4I4526_$1I4488_$1I4621_DIA[1], _4I4526_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_877_0 (_4I4526_$1I4488_$1I4621_DIA[0], _4I4526_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _4I4526_$1I4488_$1I4621_DIB;
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_878_15 (_4I4526_$1I4488_$1I4621_DIB[15], _4I4526_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_878_14 (_4I4526_$1I4488_$1I4621_DIB[14], _4I4526_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_878_13 (_4I4526_$1I4488_$1I4621_DIB[13], _4I4526_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_878_12 (_4I4526_$1I4488_$1I4621_DIB[12], _4I4526_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_878_11 (_4I4526_$1I4488_$1I4621_DIB[11], _4I4526_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_878_10 (_4I4526_$1I4488_$1I4621_DIB[10], _4I4526_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_878_9 (_4I4526_$1I4488_$1I4621_DIB[9], _4I4526_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_878_8 (_4I4526_$1I4488_$1I4621_DIB[8], _4I4526_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_878_7 (_4I4526_$1I4488_$1I4621_DIB[7], _4I4526_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_878_6 (_4I4526_$1I4488_$1I4621_DIB[6], _4I4526_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_878_5 (_4I4526_$1I4488_$1I4621_DIB[5], _4I4526_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_878_4 (_4I4526_$1I4488_$1I4621_DIB[4], _4I4526_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_878_3 (_4I4526_$1I4488_$1I4621_DIB[3], _4I4526_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_878_2 (_4I4526_$1I4488_$1I4621_DIB[2], _4I4526_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_878_1 (_4I4526_$1I4488_$1I4621_DIB[1], _4I4526_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_878_0 (_4I4526_$1I4488_$1I4621_DIB[0], _4I4526_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _4I4526_$1I4488_$1I4621_DIPA;
 reg [1:16] _4I4526_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_879_0 (_4I4526_$1I4488_$1I4621_DIPA[0], _4I4526_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _4I4526_$1I4488_$1I4621_DIPB;
 reg [1:16] _4I4526_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_880_1 (_4I4526_$1I4488_$1I4621_DIPB[1], _4I4526_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_880_0 (_4I4526_$1I4488_$1I4621_DIPB[0], _4I4526_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _4I4526_$1I4488_$1I4621_ENA;
 reg [1:16] _4I4526_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_881 (_4I4526_$1I4488_$1I4621_ENA, _4I4526_$1I4488_$1I4621_ENA__vlIN);

 wire  _4I4526_$1I4488_$1I4621_ENB;
 reg [1:16] _4I4526_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_882 (_4I4526_$1I4488_$1I4621_ENB, _4I4526_$1I4488_$1I4621_ENB__vlIN);

 wire  _4I4526_$1I4488_$1I4621_SSRA;
 reg [1:16] _4I4526_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_883 (_4I4526_$1I4488_$1I4621_SSRA, _4I4526_$1I4488_$1I4621_SSRA__vlIN);

 wire  _4I4526_$1I4488_$1I4621_SSRB;
 reg [1:16] _4I4526_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_884 (_4I4526_$1I4488_$1I4621_SSRB, _4I4526_$1I4488_$1I4621_SSRB__vlIN);

 wire  _4I4526_$1I4488_$1I4621_WEA;
 reg [1:16] _4I4526_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_885 (_4I4526_$1I4488_$1I4621_WEA, _4I4526_$1I4488_$1I4621_WEA__vlIN);

 wire  _4I4526_$1I4488_$1I4621_WEB;
 reg [1:16] _4I4526_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_886 (_4I4526_$1I4488_$1I4621_WEB, _4I4526_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _4I4526_$1I4488_$1I4621 ( _4I4526_$1I4488_$1I4621_DOA , _4I4526_$1I4488_$1I4621_DOB , _4I4526_$1I4488_$1I4621_DOPA , _4I4526_$1I4488_$1I4621_DOPB , _4I4526_$1I4488_$1I4621_ADDRA , _4I4526_$1I4488_$1I4621_ADDRB , _4I4526_$1I4488_$1I4621_CLKA , _4I4526_$1I4488_$1I4621_CLKB , _4I4526_$1I4488_$1I4621_DIA , _4I4526_$1I4488_$1I4621_DIB , _4I4526_$1I4488_$1I4621_DIPA , _4I4526_$1I4488_$1I4621_DIPB , _4I4526_$1I4488_$1I4621_ENA , _4I4526_$1I4488_$1I4621_ENB , _4I4526_$1I4488_$1I4621_SSRA , _4I4526_$1I4488_$1I4621_SSRB , _4I4526_$1I4488_$1I4621_WEA , _4I4526_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4526_$1I4488_$1I4620_DOA;

 wire [15:0] _4I4526_$1I4488_$1I4620_DOB;

 wire [0:0] _4I4526_$1I4488_$1I4620_DOPA;

 wire [1:0] _4I4526_$1I4488_$1I4620_DOPB;

 wire [10:0] _4I4526_$1I4488_$1I4620_ADDRA;
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_887_10 (_4I4526_$1I4488_$1I4620_ADDRA[10], _4I4526_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_887_9 (_4I4526_$1I4488_$1I4620_ADDRA[9], _4I4526_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_887_8 (_4I4526_$1I4488_$1I4620_ADDRA[8], _4I4526_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_887_7 (_4I4526_$1I4488_$1I4620_ADDRA[7], _4I4526_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_887_6 (_4I4526_$1I4488_$1I4620_ADDRA[6], _4I4526_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_887_5 (_4I4526_$1I4488_$1I4620_ADDRA[5], _4I4526_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_887_4 (_4I4526_$1I4488_$1I4620_ADDRA[4], _4I4526_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_887_3 (_4I4526_$1I4488_$1I4620_ADDRA[3], _4I4526_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_887_2 (_4I4526_$1I4488_$1I4620_ADDRA[2], _4I4526_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_887_1 (_4I4526_$1I4488_$1I4620_ADDRA[1], _4I4526_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_887_0 (_4I4526_$1I4488_$1I4620_ADDRA[0], _4I4526_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _4I4526_$1I4488_$1I4620_ADDRB;
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_888_9 (_4I4526_$1I4488_$1I4620_ADDRB[9], _4I4526_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_888_8 (_4I4526_$1I4488_$1I4620_ADDRB[8], _4I4526_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_888_7 (_4I4526_$1I4488_$1I4620_ADDRB[7], _4I4526_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_888_6 (_4I4526_$1I4488_$1I4620_ADDRB[6], _4I4526_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_888_5 (_4I4526_$1I4488_$1I4620_ADDRB[5], _4I4526_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_888_4 (_4I4526_$1I4488_$1I4620_ADDRB[4], _4I4526_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_888_3 (_4I4526_$1I4488_$1I4620_ADDRB[3], _4I4526_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_888_2 (_4I4526_$1I4488_$1I4620_ADDRB[2], _4I4526_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_888_1 (_4I4526_$1I4488_$1I4620_ADDRB[1], _4I4526_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_888_0 (_4I4526_$1I4488_$1I4620_ADDRB[0], _4I4526_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _4I4526_$1I4488_$1I4620_CLKA;
 reg [1:16] _4I4526_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_889 (_4I4526_$1I4488_$1I4620_CLKA, _4I4526_$1I4488_$1I4620_CLKA__vlIN);

 wire  _4I4526_$1I4488_$1I4620_CLKB;
 reg [1:16] _4I4526_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_890 (_4I4526_$1I4488_$1I4620_CLKB, _4I4526_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _4I4526_$1I4488_$1I4620_DIA;
 reg [1:16] _4I4526_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_891_7 (_4I4526_$1I4488_$1I4620_DIA[7], _4I4526_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_891_6 (_4I4526_$1I4488_$1I4620_DIA[6], _4I4526_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_891_5 (_4I4526_$1I4488_$1I4620_DIA[5], _4I4526_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_891_4 (_4I4526_$1I4488_$1I4620_DIA[4], _4I4526_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_891_3 (_4I4526_$1I4488_$1I4620_DIA[3], _4I4526_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_891_2 (_4I4526_$1I4488_$1I4620_DIA[2], _4I4526_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_891_1 (_4I4526_$1I4488_$1I4620_DIA[1], _4I4526_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_891_0 (_4I4526_$1I4488_$1I4620_DIA[0], _4I4526_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _4I4526_$1I4488_$1I4620_DIB;
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_892_15 (_4I4526_$1I4488_$1I4620_DIB[15], _4I4526_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_892_14 (_4I4526_$1I4488_$1I4620_DIB[14], _4I4526_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_892_13 (_4I4526_$1I4488_$1I4620_DIB[13], _4I4526_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_892_12 (_4I4526_$1I4488_$1I4620_DIB[12], _4I4526_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_892_11 (_4I4526_$1I4488_$1I4620_DIB[11], _4I4526_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_892_10 (_4I4526_$1I4488_$1I4620_DIB[10], _4I4526_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_892_9 (_4I4526_$1I4488_$1I4620_DIB[9], _4I4526_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_892_8 (_4I4526_$1I4488_$1I4620_DIB[8], _4I4526_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_892_7 (_4I4526_$1I4488_$1I4620_DIB[7], _4I4526_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_892_6 (_4I4526_$1I4488_$1I4620_DIB[6], _4I4526_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_892_5 (_4I4526_$1I4488_$1I4620_DIB[5], _4I4526_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_892_4 (_4I4526_$1I4488_$1I4620_DIB[4], _4I4526_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_892_3 (_4I4526_$1I4488_$1I4620_DIB[3], _4I4526_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_892_2 (_4I4526_$1I4488_$1I4620_DIB[2], _4I4526_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_892_1 (_4I4526_$1I4488_$1I4620_DIB[1], _4I4526_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_892_0 (_4I4526_$1I4488_$1I4620_DIB[0], _4I4526_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _4I4526_$1I4488_$1I4620_DIPA;
 reg [1:16] _4I4526_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_893_0 (_4I4526_$1I4488_$1I4620_DIPA[0], _4I4526_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _4I4526_$1I4488_$1I4620_DIPB;
 reg [1:16] _4I4526_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_894_1 (_4I4526_$1I4488_$1I4620_DIPB[1], _4I4526_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _4I4526_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_894_0 (_4I4526_$1I4488_$1I4620_DIPB[0], _4I4526_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _4I4526_$1I4488_$1I4620_ENA;
 reg [1:16] _4I4526_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_895 (_4I4526_$1I4488_$1I4620_ENA, _4I4526_$1I4488_$1I4620_ENA__vlIN);

 wire  _4I4526_$1I4488_$1I4620_ENB;
 reg [1:16] _4I4526_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_896 (_4I4526_$1I4488_$1I4620_ENB, _4I4526_$1I4488_$1I4620_ENB__vlIN);

 wire  _4I4526_$1I4488_$1I4620_SSRA;
 reg [1:16] _4I4526_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_897 (_4I4526_$1I4488_$1I4620_SSRA, _4I4526_$1I4488_$1I4620_SSRA__vlIN);

 wire  _4I4526_$1I4488_$1I4620_SSRB;
 reg [1:16] _4I4526_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_898 (_4I4526_$1I4488_$1I4620_SSRB, _4I4526_$1I4488_$1I4620_SSRB__vlIN);

 wire  _4I4526_$1I4488_$1I4620_WEA;
 reg [1:16] _4I4526_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_899 (_4I4526_$1I4488_$1I4620_WEA, _4I4526_$1I4488_$1I4620_WEA__vlIN);

 wire  _4I4526_$1I4488_$1I4620_WEB;
 reg [1:16] _4I4526_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_900 (_4I4526_$1I4488_$1I4620_WEB, _4I4526_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _4I4526_$1I4488_$1I4620 ( _4I4526_$1I4488_$1I4620_DOA , _4I4526_$1I4488_$1I4620_DOB , _4I4526_$1I4488_$1I4620_DOPA , _4I4526_$1I4488_$1I4620_DOPB , _4I4526_$1I4488_$1I4620_ADDRA , _4I4526_$1I4488_$1I4620_ADDRB , _4I4526_$1I4488_$1I4620_CLKA , _4I4526_$1I4488_$1I4620_CLKB , _4I4526_$1I4488_$1I4620_DIA , _4I4526_$1I4488_$1I4620_DIB , _4I4526_$1I4488_$1I4620_DIPA , _4I4526_$1I4488_$1I4620_DIPB , _4I4526_$1I4488_$1I4620_ENA , _4I4526_$1I4488_$1I4620_ENB , _4I4526_$1I4488_$1I4620_SSRA , _4I4526_$1I4488_$1I4620_SSRB , _4I4526_$1I4488_$1I4620_WEA , _4I4526_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4501_$1I4488_$1I4621_DOA;

 wire [15:0] _4I4501_$1I4488_$1I4621_DOB;

 wire [0:0] _4I4501_$1I4488_$1I4621_DOPA;

 wire [1:0] _4I4501_$1I4488_$1I4621_DOPB;

 wire [10:0] _4I4501_$1I4488_$1I4621_ADDRA;
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_901_10 (_4I4501_$1I4488_$1I4621_ADDRA[10], _4I4501_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_901_9 (_4I4501_$1I4488_$1I4621_ADDRA[9], _4I4501_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_901_8 (_4I4501_$1I4488_$1I4621_ADDRA[8], _4I4501_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_901_7 (_4I4501_$1I4488_$1I4621_ADDRA[7], _4I4501_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_901_6 (_4I4501_$1I4488_$1I4621_ADDRA[6], _4I4501_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_901_5 (_4I4501_$1I4488_$1I4621_ADDRA[5], _4I4501_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_901_4 (_4I4501_$1I4488_$1I4621_ADDRA[4], _4I4501_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_901_3 (_4I4501_$1I4488_$1I4621_ADDRA[3], _4I4501_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_901_2 (_4I4501_$1I4488_$1I4621_ADDRA[2], _4I4501_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_901_1 (_4I4501_$1I4488_$1I4621_ADDRA[1], _4I4501_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_901_0 (_4I4501_$1I4488_$1I4621_ADDRA[0], _4I4501_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _4I4501_$1I4488_$1I4621_ADDRB;
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_902_9 (_4I4501_$1I4488_$1I4621_ADDRB[9], _4I4501_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_902_8 (_4I4501_$1I4488_$1I4621_ADDRB[8], _4I4501_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_902_7 (_4I4501_$1I4488_$1I4621_ADDRB[7], _4I4501_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_902_6 (_4I4501_$1I4488_$1I4621_ADDRB[6], _4I4501_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_902_5 (_4I4501_$1I4488_$1I4621_ADDRB[5], _4I4501_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_902_4 (_4I4501_$1I4488_$1I4621_ADDRB[4], _4I4501_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_902_3 (_4I4501_$1I4488_$1I4621_ADDRB[3], _4I4501_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_902_2 (_4I4501_$1I4488_$1I4621_ADDRB[2], _4I4501_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_902_1 (_4I4501_$1I4488_$1I4621_ADDRB[1], _4I4501_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_902_0 (_4I4501_$1I4488_$1I4621_ADDRB[0], _4I4501_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _4I4501_$1I4488_$1I4621_CLKA;
 reg [1:16] _4I4501_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_903 (_4I4501_$1I4488_$1I4621_CLKA, _4I4501_$1I4488_$1I4621_CLKA__vlIN);

 wire  _4I4501_$1I4488_$1I4621_CLKB;
 reg [1:16] _4I4501_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_904 (_4I4501_$1I4488_$1I4621_CLKB, _4I4501_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _4I4501_$1I4488_$1I4621_DIA;
 reg [1:16] _4I4501_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_905_7 (_4I4501_$1I4488_$1I4621_DIA[7], _4I4501_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_905_6 (_4I4501_$1I4488_$1I4621_DIA[6], _4I4501_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_905_5 (_4I4501_$1I4488_$1I4621_DIA[5], _4I4501_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_905_4 (_4I4501_$1I4488_$1I4621_DIA[4], _4I4501_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_905_3 (_4I4501_$1I4488_$1I4621_DIA[3], _4I4501_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_905_2 (_4I4501_$1I4488_$1I4621_DIA[2], _4I4501_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_905_1 (_4I4501_$1I4488_$1I4621_DIA[1], _4I4501_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_905_0 (_4I4501_$1I4488_$1I4621_DIA[0], _4I4501_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _4I4501_$1I4488_$1I4621_DIB;
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_906_15 (_4I4501_$1I4488_$1I4621_DIB[15], _4I4501_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_906_14 (_4I4501_$1I4488_$1I4621_DIB[14], _4I4501_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_906_13 (_4I4501_$1I4488_$1I4621_DIB[13], _4I4501_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_906_12 (_4I4501_$1I4488_$1I4621_DIB[12], _4I4501_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_906_11 (_4I4501_$1I4488_$1I4621_DIB[11], _4I4501_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_906_10 (_4I4501_$1I4488_$1I4621_DIB[10], _4I4501_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_906_9 (_4I4501_$1I4488_$1I4621_DIB[9], _4I4501_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_906_8 (_4I4501_$1I4488_$1I4621_DIB[8], _4I4501_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_906_7 (_4I4501_$1I4488_$1I4621_DIB[7], _4I4501_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_906_6 (_4I4501_$1I4488_$1I4621_DIB[6], _4I4501_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_906_5 (_4I4501_$1I4488_$1I4621_DIB[5], _4I4501_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_906_4 (_4I4501_$1I4488_$1I4621_DIB[4], _4I4501_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_906_3 (_4I4501_$1I4488_$1I4621_DIB[3], _4I4501_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_906_2 (_4I4501_$1I4488_$1I4621_DIB[2], _4I4501_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_906_1 (_4I4501_$1I4488_$1I4621_DIB[1], _4I4501_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_906_0 (_4I4501_$1I4488_$1I4621_DIB[0], _4I4501_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _4I4501_$1I4488_$1I4621_DIPA;
 reg [1:16] _4I4501_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_907_0 (_4I4501_$1I4488_$1I4621_DIPA[0], _4I4501_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _4I4501_$1I4488_$1I4621_DIPB;
 reg [1:16] _4I4501_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_908_1 (_4I4501_$1I4488_$1I4621_DIPB[1], _4I4501_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_908_0 (_4I4501_$1I4488_$1I4621_DIPB[0], _4I4501_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _4I4501_$1I4488_$1I4621_ENA;
 reg [1:16] _4I4501_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_909 (_4I4501_$1I4488_$1I4621_ENA, _4I4501_$1I4488_$1I4621_ENA__vlIN);

 wire  _4I4501_$1I4488_$1I4621_ENB;
 reg [1:16] _4I4501_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_910 (_4I4501_$1I4488_$1I4621_ENB, _4I4501_$1I4488_$1I4621_ENB__vlIN);

 wire  _4I4501_$1I4488_$1I4621_SSRA;
 reg [1:16] _4I4501_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_911 (_4I4501_$1I4488_$1I4621_SSRA, _4I4501_$1I4488_$1I4621_SSRA__vlIN);

 wire  _4I4501_$1I4488_$1I4621_SSRB;
 reg [1:16] _4I4501_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_912 (_4I4501_$1I4488_$1I4621_SSRB, _4I4501_$1I4488_$1I4621_SSRB__vlIN);

 wire  _4I4501_$1I4488_$1I4621_WEA;
 reg [1:16] _4I4501_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_913 (_4I4501_$1I4488_$1I4621_WEA, _4I4501_$1I4488_$1I4621_WEA__vlIN);

 wire  _4I4501_$1I4488_$1I4621_WEB;
 reg [1:16] _4I4501_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_914 (_4I4501_$1I4488_$1I4621_WEB, _4I4501_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _4I4501_$1I4488_$1I4621 ( _4I4501_$1I4488_$1I4621_DOA , _4I4501_$1I4488_$1I4621_DOB , _4I4501_$1I4488_$1I4621_DOPA , _4I4501_$1I4488_$1I4621_DOPB , _4I4501_$1I4488_$1I4621_ADDRA , _4I4501_$1I4488_$1I4621_ADDRB , _4I4501_$1I4488_$1I4621_CLKA , _4I4501_$1I4488_$1I4621_CLKB , _4I4501_$1I4488_$1I4621_DIA , _4I4501_$1I4488_$1I4621_DIB , _4I4501_$1I4488_$1I4621_DIPA , _4I4501_$1I4488_$1I4621_DIPB , _4I4501_$1I4488_$1I4621_ENA , _4I4501_$1I4488_$1I4621_ENB , _4I4501_$1I4488_$1I4621_SSRA , _4I4501_$1I4488_$1I4621_SSRB , _4I4501_$1I4488_$1I4621_WEA , _4I4501_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4501_$1I4488_$1I4620_DOA;

 wire [15:0] _4I4501_$1I4488_$1I4620_DOB;

 wire [0:0] _4I4501_$1I4488_$1I4620_DOPA;

 wire [1:0] _4I4501_$1I4488_$1I4620_DOPB;

 wire [10:0] _4I4501_$1I4488_$1I4620_ADDRA;
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_915_10 (_4I4501_$1I4488_$1I4620_ADDRA[10], _4I4501_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_915_9 (_4I4501_$1I4488_$1I4620_ADDRA[9], _4I4501_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_915_8 (_4I4501_$1I4488_$1I4620_ADDRA[8], _4I4501_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_915_7 (_4I4501_$1I4488_$1I4620_ADDRA[7], _4I4501_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_915_6 (_4I4501_$1I4488_$1I4620_ADDRA[6], _4I4501_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_915_5 (_4I4501_$1I4488_$1I4620_ADDRA[5], _4I4501_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_915_4 (_4I4501_$1I4488_$1I4620_ADDRA[4], _4I4501_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_915_3 (_4I4501_$1I4488_$1I4620_ADDRA[3], _4I4501_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_915_2 (_4I4501_$1I4488_$1I4620_ADDRA[2], _4I4501_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_915_1 (_4I4501_$1I4488_$1I4620_ADDRA[1], _4I4501_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_915_0 (_4I4501_$1I4488_$1I4620_ADDRA[0], _4I4501_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _4I4501_$1I4488_$1I4620_ADDRB;
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_916_9 (_4I4501_$1I4488_$1I4620_ADDRB[9], _4I4501_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_916_8 (_4I4501_$1I4488_$1I4620_ADDRB[8], _4I4501_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_916_7 (_4I4501_$1I4488_$1I4620_ADDRB[7], _4I4501_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_916_6 (_4I4501_$1I4488_$1I4620_ADDRB[6], _4I4501_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_916_5 (_4I4501_$1I4488_$1I4620_ADDRB[5], _4I4501_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_916_4 (_4I4501_$1I4488_$1I4620_ADDRB[4], _4I4501_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_916_3 (_4I4501_$1I4488_$1I4620_ADDRB[3], _4I4501_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_916_2 (_4I4501_$1I4488_$1I4620_ADDRB[2], _4I4501_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_916_1 (_4I4501_$1I4488_$1I4620_ADDRB[1], _4I4501_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_916_0 (_4I4501_$1I4488_$1I4620_ADDRB[0], _4I4501_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _4I4501_$1I4488_$1I4620_CLKA;
 reg [1:16] _4I4501_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_917 (_4I4501_$1I4488_$1I4620_CLKA, _4I4501_$1I4488_$1I4620_CLKA__vlIN);

 wire  _4I4501_$1I4488_$1I4620_CLKB;
 reg [1:16] _4I4501_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_918 (_4I4501_$1I4488_$1I4620_CLKB, _4I4501_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _4I4501_$1I4488_$1I4620_DIA;
 reg [1:16] _4I4501_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_919_7 (_4I4501_$1I4488_$1I4620_DIA[7], _4I4501_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_919_6 (_4I4501_$1I4488_$1I4620_DIA[6], _4I4501_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_919_5 (_4I4501_$1I4488_$1I4620_DIA[5], _4I4501_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_919_4 (_4I4501_$1I4488_$1I4620_DIA[4], _4I4501_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_919_3 (_4I4501_$1I4488_$1I4620_DIA[3], _4I4501_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_919_2 (_4I4501_$1I4488_$1I4620_DIA[2], _4I4501_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_919_1 (_4I4501_$1I4488_$1I4620_DIA[1], _4I4501_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_919_0 (_4I4501_$1I4488_$1I4620_DIA[0], _4I4501_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _4I4501_$1I4488_$1I4620_DIB;
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_920_15 (_4I4501_$1I4488_$1I4620_DIB[15], _4I4501_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_920_14 (_4I4501_$1I4488_$1I4620_DIB[14], _4I4501_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_920_13 (_4I4501_$1I4488_$1I4620_DIB[13], _4I4501_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_920_12 (_4I4501_$1I4488_$1I4620_DIB[12], _4I4501_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_920_11 (_4I4501_$1I4488_$1I4620_DIB[11], _4I4501_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_920_10 (_4I4501_$1I4488_$1I4620_DIB[10], _4I4501_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_920_9 (_4I4501_$1I4488_$1I4620_DIB[9], _4I4501_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_920_8 (_4I4501_$1I4488_$1I4620_DIB[8], _4I4501_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_920_7 (_4I4501_$1I4488_$1I4620_DIB[7], _4I4501_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_920_6 (_4I4501_$1I4488_$1I4620_DIB[6], _4I4501_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_920_5 (_4I4501_$1I4488_$1I4620_DIB[5], _4I4501_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_920_4 (_4I4501_$1I4488_$1I4620_DIB[4], _4I4501_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_920_3 (_4I4501_$1I4488_$1I4620_DIB[3], _4I4501_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_920_2 (_4I4501_$1I4488_$1I4620_DIB[2], _4I4501_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_920_1 (_4I4501_$1I4488_$1I4620_DIB[1], _4I4501_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_920_0 (_4I4501_$1I4488_$1I4620_DIB[0], _4I4501_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _4I4501_$1I4488_$1I4620_DIPA;
 reg [1:16] _4I4501_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_921_0 (_4I4501_$1I4488_$1I4620_DIPA[0], _4I4501_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _4I4501_$1I4488_$1I4620_DIPB;
 reg [1:16] _4I4501_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_922_1 (_4I4501_$1I4488_$1I4620_DIPB[1], _4I4501_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _4I4501_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_922_0 (_4I4501_$1I4488_$1I4620_DIPB[0], _4I4501_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _4I4501_$1I4488_$1I4620_ENA;
 reg [1:16] _4I4501_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_923 (_4I4501_$1I4488_$1I4620_ENA, _4I4501_$1I4488_$1I4620_ENA__vlIN);

 wire  _4I4501_$1I4488_$1I4620_ENB;
 reg [1:16] _4I4501_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_924 (_4I4501_$1I4488_$1I4620_ENB, _4I4501_$1I4488_$1I4620_ENB__vlIN);

 wire  _4I4501_$1I4488_$1I4620_SSRA;
 reg [1:16] _4I4501_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_925 (_4I4501_$1I4488_$1I4620_SSRA, _4I4501_$1I4488_$1I4620_SSRA__vlIN);

 wire  _4I4501_$1I4488_$1I4620_SSRB;
 reg [1:16] _4I4501_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_926 (_4I4501_$1I4488_$1I4620_SSRB, _4I4501_$1I4488_$1I4620_SSRB__vlIN);

 wire  _4I4501_$1I4488_$1I4620_WEA;
 reg [1:16] _4I4501_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_927 (_4I4501_$1I4488_$1I4620_WEA, _4I4501_$1I4488_$1I4620_WEA__vlIN);

 wire  _4I4501_$1I4488_$1I4620_WEB;
 reg [1:16] _4I4501_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_928 (_4I4501_$1I4488_$1I4620_WEB, _4I4501_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _4I4501_$1I4488_$1I4620 ( _4I4501_$1I4488_$1I4620_DOA , _4I4501_$1I4488_$1I4620_DOB , _4I4501_$1I4488_$1I4620_DOPA , _4I4501_$1I4488_$1I4620_DOPB , _4I4501_$1I4488_$1I4620_ADDRA , _4I4501_$1I4488_$1I4620_ADDRB , _4I4501_$1I4488_$1I4620_CLKA , _4I4501_$1I4488_$1I4620_CLKB , _4I4501_$1I4488_$1I4620_DIA , _4I4501_$1I4488_$1I4620_DIB , _4I4501_$1I4488_$1I4620_DIPA , _4I4501_$1I4488_$1I4620_DIPB , _4I4501_$1I4488_$1I4620_ENA , _4I4501_$1I4488_$1I4620_ENB , _4I4501_$1I4488_$1I4620_SSRA , _4I4501_$1I4488_$1I4620_SSRB , _4I4501_$1I4488_$1I4620_WEA , _4I4501_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4476_$1I4488_$1I4621_DOA;

 wire [15:0] _4I4476_$1I4488_$1I4621_DOB;

 wire [0:0] _4I4476_$1I4488_$1I4621_DOPA;

 wire [1:0] _4I4476_$1I4488_$1I4621_DOPB;

 wire [10:0] _4I4476_$1I4488_$1I4621_ADDRA;
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_929_10 (_4I4476_$1I4488_$1I4621_ADDRA[10], _4I4476_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_929_9 (_4I4476_$1I4488_$1I4621_ADDRA[9], _4I4476_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_929_8 (_4I4476_$1I4488_$1I4621_ADDRA[8], _4I4476_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_929_7 (_4I4476_$1I4488_$1I4621_ADDRA[7], _4I4476_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_929_6 (_4I4476_$1I4488_$1I4621_ADDRA[6], _4I4476_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_929_5 (_4I4476_$1I4488_$1I4621_ADDRA[5], _4I4476_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_929_4 (_4I4476_$1I4488_$1I4621_ADDRA[4], _4I4476_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_929_3 (_4I4476_$1I4488_$1I4621_ADDRA[3], _4I4476_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_929_2 (_4I4476_$1I4488_$1I4621_ADDRA[2], _4I4476_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_929_1 (_4I4476_$1I4488_$1I4621_ADDRA[1], _4I4476_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_929_0 (_4I4476_$1I4488_$1I4621_ADDRA[0], _4I4476_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _4I4476_$1I4488_$1I4621_ADDRB;
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_930_9 (_4I4476_$1I4488_$1I4621_ADDRB[9], _4I4476_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_930_8 (_4I4476_$1I4488_$1I4621_ADDRB[8], _4I4476_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_930_7 (_4I4476_$1I4488_$1I4621_ADDRB[7], _4I4476_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_930_6 (_4I4476_$1I4488_$1I4621_ADDRB[6], _4I4476_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_930_5 (_4I4476_$1I4488_$1I4621_ADDRB[5], _4I4476_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_930_4 (_4I4476_$1I4488_$1I4621_ADDRB[4], _4I4476_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_930_3 (_4I4476_$1I4488_$1I4621_ADDRB[3], _4I4476_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_930_2 (_4I4476_$1I4488_$1I4621_ADDRB[2], _4I4476_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_930_1 (_4I4476_$1I4488_$1I4621_ADDRB[1], _4I4476_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_930_0 (_4I4476_$1I4488_$1I4621_ADDRB[0], _4I4476_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _4I4476_$1I4488_$1I4621_CLKA;
 reg [1:16] _4I4476_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_931 (_4I4476_$1I4488_$1I4621_CLKA, _4I4476_$1I4488_$1I4621_CLKA__vlIN);

 wire  _4I4476_$1I4488_$1I4621_CLKB;
 reg [1:16] _4I4476_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_932 (_4I4476_$1I4488_$1I4621_CLKB, _4I4476_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _4I4476_$1I4488_$1I4621_DIA;
 reg [1:16] _4I4476_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_933_7 (_4I4476_$1I4488_$1I4621_DIA[7], _4I4476_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_933_6 (_4I4476_$1I4488_$1I4621_DIA[6], _4I4476_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_933_5 (_4I4476_$1I4488_$1I4621_DIA[5], _4I4476_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_933_4 (_4I4476_$1I4488_$1I4621_DIA[4], _4I4476_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_933_3 (_4I4476_$1I4488_$1I4621_DIA[3], _4I4476_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_933_2 (_4I4476_$1I4488_$1I4621_DIA[2], _4I4476_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_933_1 (_4I4476_$1I4488_$1I4621_DIA[1], _4I4476_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_933_0 (_4I4476_$1I4488_$1I4621_DIA[0], _4I4476_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _4I4476_$1I4488_$1I4621_DIB;
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_934_15 (_4I4476_$1I4488_$1I4621_DIB[15], _4I4476_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_934_14 (_4I4476_$1I4488_$1I4621_DIB[14], _4I4476_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_934_13 (_4I4476_$1I4488_$1I4621_DIB[13], _4I4476_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_934_12 (_4I4476_$1I4488_$1I4621_DIB[12], _4I4476_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_934_11 (_4I4476_$1I4488_$1I4621_DIB[11], _4I4476_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_934_10 (_4I4476_$1I4488_$1I4621_DIB[10], _4I4476_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_934_9 (_4I4476_$1I4488_$1I4621_DIB[9], _4I4476_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_934_8 (_4I4476_$1I4488_$1I4621_DIB[8], _4I4476_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_934_7 (_4I4476_$1I4488_$1I4621_DIB[7], _4I4476_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_934_6 (_4I4476_$1I4488_$1I4621_DIB[6], _4I4476_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_934_5 (_4I4476_$1I4488_$1I4621_DIB[5], _4I4476_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_934_4 (_4I4476_$1I4488_$1I4621_DIB[4], _4I4476_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_934_3 (_4I4476_$1I4488_$1I4621_DIB[3], _4I4476_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_934_2 (_4I4476_$1I4488_$1I4621_DIB[2], _4I4476_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_934_1 (_4I4476_$1I4488_$1I4621_DIB[1], _4I4476_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_934_0 (_4I4476_$1I4488_$1I4621_DIB[0], _4I4476_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _4I4476_$1I4488_$1I4621_DIPA;
 reg [1:16] _4I4476_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_935_0 (_4I4476_$1I4488_$1I4621_DIPA[0], _4I4476_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _4I4476_$1I4488_$1I4621_DIPB;
 reg [1:16] _4I4476_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_936_1 (_4I4476_$1I4488_$1I4621_DIPB[1], _4I4476_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_936_0 (_4I4476_$1I4488_$1I4621_DIPB[0], _4I4476_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _4I4476_$1I4488_$1I4621_ENA;
 reg [1:16] _4I4476_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_937 (_4I4476_$1I4488_$1I4621_ENA, _4I4476_$1I4488_$1I4621_ENA__vlIN);

 wire  _4I4476_$1I4488_$1I4621_ENB;
 reg [1:16] _4I4476_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_938 (_4I4476_$1I4488_$1I4621_ENB, _4I4476_$1I4488_$1I4621_ENB__vlIN);

 wire  _4I4476_$1I4488_$1I4621_SSRA;
 reg [1:16] _4I4476_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_939 (_4I4476_$1I4488_$1I4621_SSRA, _4I4476_$1I4488_$1I4621_SSRA__vlIN);

 wire  _4I4476_$1I4488_$1I4621_SSRB;
 reg [1:16] _4I4476_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_940 (_4I4476_$1I4488_$1I4621_SSRB, _4I4476_$1I4488_$1I4621_SSRB__vlIN);

 wire  _4I4476_$1I4488_$1I4621_WEA;
 reg [1:16] _4I4476_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_941 (_4I4476_$1I4488_$1I4621_WEA, _4I4476_$1I4488_$1I4621_WEA__vlIN);

 wire  _4I4476_$1I4488_$1I4621_WEB;
 reg [1:16] _4I4476_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_942 (_4I4476_$1I4488_$1I4621_WEB, _4I4476_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _4I4476_$1I4488_$1I4621 ( _4I4476_$1I4488_$1I4621_DOA , _4I4476_$1I4488_$1I4621_DOB , _4I4476_$1I4488_$1I4621_DOPA , _4I4476_$1I4488_$1I4621_DOPB , _4I4476_$1I4488_$1I4621_ADDRA , _4I4476_$1I4488_$1I4621_ADDRB , _4I4476_$1I4488_$1I4621_CLKA , _4I4476_$1I4488_$1I4621_CLKB , _4I4476_$1I4488_$1I4621_DIA , _4I4476_$1I4488_$1I4621_DIB , _4I4476_$1I4488_$1I4621_DIPA , _4I4476_$1I4488_$1I4621_DIPB , _4I4476_$1I4488_$1I4621_ENA , _4I4476_$1I4488_$1I4621_ENB , _4I4476_$1I4488_$1I4621_SSRA , _4I4476_$1I4488_$1I4621_SSRB , _4I4476_$1I4488_$1I4621_WEA , _4I4476_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4476_$1I4488_$1I4620_DOA;

 wire [15:0] _4I4476_$1I4488_$1I4620_DOB;

 wire [0:0] _4I4476_$1I4488_$1I4620_DOPA;

 wire [1:0] _4I4476_$1I4488_$1I4620_DOPB;

 wire [10:0] _4I4476_$1I4488_$1I4620_ADDRA;
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_943_10 (_4I4476_$1I4488_$1I4620_ADDRA[10], _4I4476_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_943_9 (_4I4476_$1I4488_$1I4620_ADDRA[9], _4I4476_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_943_8 (_4I4476_$1I4488_$1I4620_ADDRA[8], _4I4476_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_943_7 (_4I4476_$1I4488_$1I4620_ADDRA[7], _4I4476_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_943_6 (_4I4476_$1I4488_$1I4620_ADDRA[6], _4I4476_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_943_5 (_4I4476_$1I4488_$1I4620_ADDRA[5], _4I4476_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_943_4 (_4I4476_$1I4488_$1I4620_ADDRA[4], _4I4476_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_943_3 (_4I4476_$1I4488_$1I4620_ADDRA[3], _4I4476_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_943_2 (_4I4476_$1I4488_$1I4620_ADDRA[2], _4I4476_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_943_1 (_4I4476_$1I4488_$1I4620_ADDRA[1], _4I4476_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_943_0 (_4I4476_$1I4488_$1I4620_ADDRA[0], _4I4476_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _4I4476_$1I4488_$1I4620_ADDRB;
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_944_9 (_4I4476_$1I4488_$1I4620_ADDRB[9], _4I4476_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_944_8 (_4I4476_$1I4488_$1I4620_ADDRB[8], _4I4476_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_944_7 (_4I4476_$1I4488_$1I4620_ADDRB[7], _4I4476_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_944_6 (_4I4476_$1I4488_$1I4620_ADDRB[6], _4I4476_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_944_5 (_4I4476_$1I4488_$1I4620_ADDRB[5], _4I4476_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_944_4 (_4I4476_$1I4488_$1I4620_ADDRB[4], _4I4476_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_944_3 (_4I4476_$1I4488_$1I4620_ADDRB[3], _4I4476_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_944_2 (_4I4476_$1I4488_$1I4620_ADDRB[2], _4I4476_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_944_1 (_4I4476_$1I4488_$1I4620_ADDRB[1], _4I4476_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_944_0 (_4I4476_$1I4488_$1I4620_ADDRB[0], _4I4476_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _4I4476_$1I4488_$1I4620_CLKA;
 reg [1:16] _4I4476_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_945 (_4I4476_$1I4488_$1I4620_CLKA, _4I4476_$1I4488_$1I4620_CLKA__vlIN);

 wire  _4I4476_$1I4488_$1I4620_CLKB;
 reg [1:16] _4I4476_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_946 (_4I4476_$1I4488_$1I4620_CLKB, _4I4476_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _4I4476_$1I4488_$1I4620_DIA;
 reg [1:16] _4I4476_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_947_7 (_4I4476_$1I4488_$1I4620_DIA[7], _4I4476_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_947_6 (_4I4476_$1I4488_$1I4620_DIA[6], _4I4476_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_947_5 (_4I4476_$1I4488_$1I4620_DIA[5], _4I4476_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_947_4 (_4I4476_$1I4488_$1I4620_DIA[4], _4I4476_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_947_3 (_4I4476_$1I4488_$1I4620_DIA[3], _4I4476_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_947_2 (_4I4476_$1I4488_$1I4620_DIA[2], _4I4476_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_947_1 (_4I4476_$1I4488_$1I4620_DIA[1], _4I4476_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_947_0 (_4I4476_$1I4488_$1I4620_DIA[0], _4I4476_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _4I4476_$1I4488_$1I4620_DIB;
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_948_15 (_4I4476_$1I4488_$1I4620_DIB[15], _4I4476_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_948_14 (_4I4476_$1I4488_$1I4620_DIB[14], _4I4476_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_948_13 (_4I4476_$1I4488_$1I4620_DIB[13], _4I4476_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_948_12 (_4I4476_$1I4488_$1I4620_DIB[12], _4I4476_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_948_11 (_4I4476_$1I4488_$1I4620_DIB[11], _4I4476_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_948_10 (_4I4476_$1I4488_$1I4620_DIB[10], _4I4476_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_948_9 (_4I4476_$1I4488_$1I4620_DIB[9], _4I4476_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_948_8 (_4I4476_$1I4488_$1I4620_DIB[8], _4I4476_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_948_7 (_4I4476_$1I4488_$1I4620_DIB[7], _4I4476_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_948_6 (_4I4476_$1I4488_$1I4620_DIB[6], _4I4476_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_948_5 (_4I4476_$1I4488_$1I4620_DIB[5], _4I4476_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_948_4 (_4I4476_$1I4488_$1I4620_DIB[4], _4I4476_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_948_3 (_4I4476_$1I4488_$1I4620_DIB[3], _4I4476_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_948_2 (_4I4476_$1I4488_$1I4620_DIB[2], _4I4476_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_948_1 (_4I4476_$1I4488_$1I4620_DIB[1], _4I4476_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_948_0 (_4I4476_$1I4488_$1I4620_DIB[0], _4I4476_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _4I4476_$1I4488_$1I4620_DIPA;
 reg [1:16] _4I4476_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_949_0 (_4I4476_$1I4488_$1I4620_DIPA[0], _4I4476_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _4I4476_$1I4488_$1I4620_DIPB;
 reg [1:16] _4I4476_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_950_1 (_4I4476_$1I4488_$1I4620_DIPB[1], _4I4476_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _4I4476_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_950_0 (_4I4476_$1I4488_$1I4620_DIPB[0], _4I4476_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _4I4476_$1I4488_$1I4620_ENA;
 reg [1:16] _4I4476_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_951 (_4I4476_$1I4488_$1I4620_ENA, _4I4476_$1I4488_$1I4620_ENA__vlIN);

 wire  _4I4476_$1I4488_$1I4620_ENB;
 reg [1:16] _4I4476_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_952 (_4I4476_$1I4488_$1I4620_ENB, _4I4476_$1I4488_$1I4620_ENB__vlIN);

 wire  _4I4476_$1I4488_$1I4620_SSRA;
 reg [1:16] _4I4476_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_953 (_4I4476_$1I4488_$1I4620_SSRA, _4I4476_$1I4488_$1I4620_SSRA__vlIN);

 wire  _4I4476_$1I4488_$1I4620_SSRB;
 reg [1:16] _4I4476_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_954 (_4I4476_$1I4488_$1I4620_SSRB, _4I4476_$1I4488_$1I4620_SSRB__vlIN);

 wire  _4I4476_$1I4488_$1I4620_WEA;
 reg [1:16] _4I4476_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_955 (_4I4476_$1I4488_$1I4620_WEA, _4I4476_$1I4488_$1I4620_WEA__vlIN);

 wire  _4I4476_$1I4488_$1I4620_WEB;
 reg [1:16] _4I4476_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_956 (_4I4476_$1I4488_$1I4620_WEB, _4I4476_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _4I4476_$1I4488_$1I4620 ( _4I4476_$1I4488_$1I4620_DOA , _4I4476_$1I4488_$1I4620_DOB , _4I4476_$1I4488_$1I4620_DOPA , _4I4476_$1I4488_$1I4620_DOPB , _4I4476_$1I4488_$1I4620_ADDRA , _4I4476_$1I4488_$1I4620_ADDRB , _4I4476_$1I4488_$1I4620_CLKA , _4I4476_$1I4488_$1I4620_CLKB , _4I4476_$1I4488_$1I4620_DIA , _4I4476_$1I4488_$1I4620_DIB , _4I4476_$1I4488_$1I4620_DIPA , _4I4476_$1I4488_$1I4620_DIPB , _4I4476_$1I4488_$1I4620_ENA , _4I4476_$1I4488_$1I4620_ENB , _4I4476_$1I4488_$1I4620_SSRA , _4I4476_$1I4488_$1I4620_SSRB , _4I4476_$1I4488_$1I4620_WEA , _4I4476_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4475_$1I4488_$1I4621_DOA;

 wire [15:0] _4I4475_$1I4488_$1I4621_DOB;

 wire [0:0] _4I4475_$1I4488_$1I4621_DOPA;

 wire [1:0] _4I4475_$1I4488_$1I4621_DOPB;

 wire [10:0] _4I4475_$1I4488_$1I4621_ADDRA;
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_957_10 (_4I4475_$1I4488_$1I4621_ADDRA[10], _4I4475_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_957_9 (_4I4475_$1I4488_$1I4621_ADDRA[9], _4I4475_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_957_8 (_4I4475_$1I4488_$1I4621_ADDRA[8], _4I4475_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_957_7 (_4I4475_$1I4488_$1I4621_ADDRA[7], _4I4475_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_957_6 (_4I4475_$1I4488_$1I4621_ADDRA[6], _4I4475_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_957_5 (_4I4475_$1I4488_$1I4621_ADDRA[5], _4I4475_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_957_4 (_4I4475_$1I4488_$1I4621_ADDRA[4], _4I4475_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_957_3 (_4I4475_$1I4488_$1I4621_ADDRA[3], _4I4475_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_957_2 (_4I4475_$1I4488_$1I4621_ADDRA[2], _4I4475_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_957_1 (_4I4475_$1I4488_$1I4621_ADDRA[1], _4I4475_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_957_0 (_4I4475_$1I4488_$1I4621_ADDRA[0], _4I4475_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _4I4475_$1I4488_$1I4621_ADDRB;
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_958_9 (_4I4475_$1I4488_$1I4621_ADDRB[9], _4I4475_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_958_8 (_4I4475_$1I4488_$1I4621_ADDRB[8], _4I4475_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_958_7 (_4I4475_$1I4488_$1I4621_ADDRB[7], _4I4475_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_958_6 (_4I4475_$1I4488_$1I4621_ADDRB[6], _4I4475_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_958_5 (_4I4475_$1I4488_$1I4621_ADDRB[5], _4I4475_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_958_4 (_4I4475_$1I4488_$1I4621_ADDRB[4], _4I4475_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_958_3 (_4I4475_$1I4488_$1I4621_ADDRB[3], _4I4475_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_958_2 (_4I4475_$1I4488_$1I4621_ADDRB[2], _4I4475_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_958_1 (_4I4475_$1I4488_$1I4621_ADDRB[1], _4I4475_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_958_0 (_4I4475_$1I4488_$1I4621_ADDRB[0], _4I4475_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _4I4475_$1I4488_$1I4621_CLKA;
 reg [1:16] _4I4475_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_959 (_4I4475_$1I4488_$1I4621_CLKA, _4I4475_$1I4488_$1I4621_CLKA__vlIN);

 wire  _4I4475_$1I4488_$1I4621_CLKB;
 reg [1:16] _4I4475_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_960 (_4I4475_$1I4488_$1I4621_CLKB, _4I4475_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _4I4475_$1I4488_$1I4621_DIA;
 reg [1:16] _4I4475_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_961_7 (_4I4475_$1I4488_$1I4621_DIA[7], _4I4475_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_961_6 (_4I4475_$1I4488_$1I4621_DIA[6], _4I4475_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_961_5 (_4I4475_$1I4488_$1I4621_DIA[5], _4I4475_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_961_4 (_4I4475_$1I4488_$1I4621_DIA[4], _4I4475_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_961_3 (_4I4475_$1I4488_$1I4621_DIA[3], _4I4475_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_961_2 (_4I4475_$1I4488_$1I4621_DIA[2], _4I4475_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_961_1 (_4I4475_$1I4488_$1I4621_DIA[1], _4I4475_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_961_0 (_4I4475_$1I4488_$1I4621_DIA[0], _4I4475_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _4I4475_$1I4488_$1I4621_DIB;
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_962_15 (_4I4475_$1I4488_$1I4621_DIB[15], _4I4475_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_962_14 (_4I4475_$1I4488_$1I4621_DIB[14], _4I4475_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_962_13 (_4I4475_$1I4488_$1I4621_DIB[13], _4I4475_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_962_12 (_4I4475_$1I4488_$1I4621_DIB[12], _4I4475_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_962_11 (_4I4475_$1I4488_$1I4621_DIB[11], _4I4475_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_962_10 (_4I4475_$1I4488_$1I4621_DIB[10], _4I4475_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_962_9 (_4I4475_$1I4488_$1I4621_DIB[9], _4I4475_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_962_8 (_4I4475_$1I4488_$1I4621_DIB[8], _4I4475_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_962_7 (_4I4475_$1I4488_$1I4621_DIB[7], _4I4475_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_962_6 (_4I4475_$1I4488_$1I4621_DIB[6], _4I4475_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_962_5 (_4I4475_$1I4488_$1I4621_DIB[5], _4I4475_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_962_4 (_4I4475_$1I4488_$1I4621_DIB[4], _4I4475_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_962_3 (_4I4475_$1I4488_$1I4621_DIB[3], _4I4475_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_962_2 (_4I4475_$1I4488_$1I4621_DIB[2], _4I4475_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_962_1 (_4I4475_$1I4488_$1I4621_DIB[1], _4I4475_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_962_0 (_4I4475_$1I4488_$1I4621_DIB[0], _4I4475_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _4I4475_$1I4488_$1I4621_DIPA;
 reg [1:16] _4I4475_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_963_0 (_4I4475_$1I4488_$1I4621_DIPA[0], _4I4475_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _4I4475_$1I4488_$1I4621_DIPB;
 reg [1:16] _4I4475_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_964_1 (_4I4475_$1I4488_$1I4621_DIPB[1], _4I4475_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_964_0 (_4I4475_$1I4488_$1I4621_DIPB[0], _4I4475_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _4I4475_$1I4488_$1I4621_ENA;
 reg [1:16] _4I4475_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_965 (_4I4475_$1I4488_$1I4621_ENA, _4I4475_$1I4488_$1I4621_ENA__vlIN);

 wire  _4I4475_$1I4488_$1I4621_ENB;
 reg [1:16] _4I4475_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_966 (_4I4475_$1I4488_$1I4621_ENB, _4I4475_$1I4488_$1I4621_ENB__vlIN);

 wire  _4I4475_$1I4488_$1I4621_SSRA;
 reg [1:16] _4I4475_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_967 (_4I4475_$1I4488_$1I4621_SSRA, _4I4475_$1I4488_$1I4621_SSRA__vlIN);

 wire  _4I4475_$1I4488_$1I4621_SSRB;
 reg [1:16] _4I4475_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_968 (_4I4475_$1I4488_$1I4621_SSRB, _4I4475_$1I4488_$1I4621_SSRB__vlIN);

 wire  _4I4475_$1I4488_$1I4621_WEA;
 reg [1:16] _4I4475_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_969 (_4I4475_$1I4488_$1I4621_WEA, _4I4475_$1I4488_$1I4621_WEA__vlIN);

 wire  _4I4475_$1I4488_$1I4621_WEB;
 reg [1:16] _4I4475_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_970 (_4I4475_$1I4488_$1I4621_WEB, _4I4475_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _4I4475_$1I4488_$1I4621 ( _4I4475_$1I4488_$1I4621_DOA , _4I4475_$1I4488_$1I4621_DOB , _4I4475_$1I4488_$1I4621_DOPA , _4I4475_$1I4488_$1I4621_DOPB , _4I4475_$1I4488_$1I4621_ADDRA , _4I4475_$1I4488_$1I4621_ADDRB , _4I4475_$1I4488_$1I4621_CLKA , _4I4475_$1I4488_$1I4621_CLKB , _4I4475_$1I4488_$1I4621_DIA , _4I4475_$1I4488_$1I4621_DIB , _4I4475_$1I4488_$1I4621_DIPA , _4I4475_$1I4488_$1I4621_DIPB , _4I4475_$1I4488_$1I4621_ENA , _4I4475_$1I4488_$1I4621_ENB , _4I4475_$1I4488_$1I4621_SSRA , _4I4475_$1I4488_$1I4621_SSRB , _4I4475_$1I4488_$1I4621_WEA , _4I4475_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4475_$1I4488_$1I4620_DOA;

 wire [15:0] _4I4475_$1I4488_$1I4620_DOB;

 wire [0:0] _4I4475_$1I4488_$1I4620_DOPA;

 wire [1:0] _4I4475_$1I4488_$1I4620_DOPB;

 wire [10:0] _4I4475_$1I4488_$1I4620_ADDRA;
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_971_10 (_4I4475_$1I4488_$1I4620_ADDRA[10], _4I4475_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_971_9 (_4I4475_$1I4488_$1I4620_ADDRA[9], _4I4475_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_971_8 (_4I4475_$1I4488_$1I4620_ADDRA[8], _4I4475_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_971_7 (_4I4475_$1I4488_$1I4620_ADDRA[7], _4I4475_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_971_6 (_4I4475_$1I4488_$1I4620_ADDRA[6], _4I4475_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_971_5 (_4I4475_$1I4488_$1I4620_ADDRA[5], _4I4475_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_971_4 (_4I4475_$1I4488_$1I4620_ADDRA[4], _4I4475_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_971_3 (_4I4475_$1I4488_$1I4620_ADDRA[3], _4I4475_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_971_2 (_4I4475_$1I4488_$1I4620_ADDRA[2], _4I4475_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_971_1 (_4I4475_$1I4488_$1I4620_ADDRA[1], _4I4475_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_971_0 (_4I4475_$1I4488_$1I4620_ADDRA[0], _4I4475_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _4I4475_$1I4488_$1I4620_ADDRB;
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_972_9 (_4I4475_$1I4488_$1I4620_ADDRB[9], _4I4475_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_972_8 (_4I4475_$1I4488_$1I4620_ADDRB[8], _4I4475_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_972_7 (_4I4475_$1I4488_$1I4620_ADDRB[7], _4I4475_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_972_6 (_4I4475_$1I4488_$1I4620_ADDRB[6], _4I4475_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_972_5 (_4I4475_$1I4488_$1I4620_ADDRB[5], _4I4475_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_972_4 (_4I4475_$1I4488_$1I4620_ADDRB[4], _4I4475_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_972_3 (_4I4475_$1I4488_$1I4620_ADDRB[3], _4I4475_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_972_2 (_4I4475_$1I4488_$1I4620_ADDRB[2], _4I4475_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_972_1 (_4I4475_$1I4488_$1I4620_ADDRB[1], _4I4475_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_972_0 (_4I4475_$1I4488_$1I4620_ADDRB[0], _4I4475_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _4I4475_$1I4488_$1I4620_CLKA;
 reg [1:16] _4I4475_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_973 (_4I4475_$1I4488_$1I4620_CLKA, _4I4475_$1I4488_$1I4620_CLKA__vlIN);

 wire  _4I4475_$1I4488_$1I4620_CLKB;
 reg [1:16] _4I4475_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_974 (_4I4475_$1I4488_$1I4620_CLKB, _4I4475_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _4I4475_$1I4488_$1I4620_DIA;
 reg [1:16] _4I4475_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_975_7 (_4I4475_$1I4488_$1I4620_DIA[7], _4I4475_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_975_6 (_4I4475_$1I4488_$1I4620_DIA[6], _4I4475_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_975_5 (_4I4475_$1I4488_$1I4620_DIA[5], _4I4475_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_975_4 (_4I4475_$1I4488_$1I4620_DIA[4], _4I4475_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_975_3 (_4I4475_$1I4488_$1I4620_DIA[3], _4I4475_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_975_2 (_4I4475_$1I4488_$1I4620_DIA[2], _4I4475_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_975_1 (_4I4475_$1I4488_$1I4620_DIA[1], _4I4475_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_975_0 (_4I4475_$1I4488_$1I4620_DIA[0], _4I4475_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _4I4475_$1I4488_$1I4620_DIB;
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_976_15 (_4I4475_$1I4488_$1I4620_DIB[15], _4I4475_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_976_14 (_4I4475_$1I4488_$1I4620_DIB[14], _4I4475_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_976_13 (_4I4475_$1I4488_$1I4620_DIB[13], _4I4475_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_976_12 (_4I4475_$1I4488_$1I4620_DIB[12], _4I4475_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_976_11 (_4I4475_$1I4488_$1I4620_DIB[11], _4I4475_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_976_10 (_4I4475_$1I4488_$1I4620_DIB[10], _4I4475_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_976_9 (_4I4475_$1I4488_$1I4620_DIB[9], _4I4475_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_976_8 (_4I4475_$1I4488_$1I4620_DIB[8], _4I4475_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_976_7 (_4I4475_$1I4488_$1I4620_DIB[7], _4I4475_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_976_6 (_4I4475_$1I4488_$1I4620_DIB[6], _4I4475_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_976_5 (_4I4475_$1I4488_$1I4620_DIB[5], _4I4475_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_976_4 (_4I4475_$1I4488_$1I4620_DIB[4], _4I4475_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_976_3 (_4I4475_$1I4488_$1I4620_DIB[3], _4I4475_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_976_2 (_4I4475_$1I4488_$1I4620_DIB[2], _4I4475_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_976_1 (_4I4475_$1I4488_$1I4620_DIB[1], _4I4475_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_976_0 (_4I4475_$1I4488_$1I4620_DIB[0], _4I4475_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _4I4475_$1I4488_$1I4620_DIPA;
 reg [1:16] _4I4475_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_977_0 (_4I4475_$1I4488_$1I4620_DIPA[0], _4I4475_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _4I4475_$1I4488_$1I4620_DIPB;
 reg [1:16] _4I4475_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_978_1 (_4I4475_$1I4488_$1I4620_DIPB[1], _4I4475_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _4I4475_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_978_0 (_4I4475_$1I4488_$1I4620_DIPB[0], _4I4475_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _4I4475_$1I4488_$1I4620_ENA;
 reg [1:16] _4I4475_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_979 (_4I4475_$1I4488_$1I4620_ENA, _4I4475_$1I4488_$1I4620_ENA__vlIN);

 wire  _4I4475_$1I4488_$1I4620_ENB;
 reg [1:16] _4I4475_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_980 (_4I4475_$1I4488_$1I4620_ENB, _4I4475_$1I4488_$1I4620_ENB__vlIN);

 wire  _4I4475_$1I4488_$1I4620_SSRA;
 reg [1:16] _4I4475_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_981 (_4I4475_$1I4488_$1I4620_SSRA, _4I4475_$1I4488_$1I4620_SSRA__vlIN);

 wire  _4I4475_$1I4488_$1I4620_SSRB;
 reg [1:16] _4I4475_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_982 (_4I4475_$1I4488_$1I4620_SSRB, _4I4475_$1I4488_$1I4620_SSRB__vlIN);

 wire  _4I4475_$1I4488_$1I4620_WEA;
 reg [1:16] _4I4475_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_983 (_4I4475_$1I4488_$1I4620_WEA, _4I4475_$1I4488_$1I4620_WEA__vlIN);

 wire  _4I4475_$1I4488_$1I4620_WEB;
 reg [1:16] _4I4475_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_984 (_4I4475_$1I4488_$1I4620_WEB, _4I4475_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _4I4475_$1I4488_$1I4620 ( _4I4475_$1I4488_$1I4620_DOA , _4I4475_$1I4488_$1I4620_DOB , _4I4475_$1I4488_$1I4620_DOPA , _4I4475_$1I4488_$1I4620_DOPB , _4I4475_$1I4488_$1I4620_ADDRA , _4I4475_$1I4488_$1I4620_ADDRB , _4I4475_$1I4488_$1I4620_CLKA , _4I4475_$1I4488_$1I4620_CLKB , _4I4475_$1I4488_$1I4620_DIA , _4I4475_$1I4488_$1I4620_DIB , _4I4475_$1I4488_$1I4620_DIPA , _4I4475_$1I4488_$1I4620_DIPB , _4I4475_$1I4488_$1I4620_ENA , _4I4475_$1I4488_$1I4620_ENB , _4I4475_$1I4488_$1I4620_SSRA , _4I4475_$1I4488_$1I4620_SSRB , _4I4475_$1I4488_$1I4620_WEA , _4I4475_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4426_$1I4488_$1I4621_DOA;

 wire [15:0] _4I4426_$1I4488_$1I4621_DOB;

 wire [0:0] _4I4426_$1I4488_$1I4621_DOPA;

 wire [1:0] _4I4426_$1I4488_$1I4621_DOPB;

 wire [10:0] _4I4426_$1I4488_$1I4621_ADDRA;
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_985_10 (_4I4426_$1I4488_$1I4621_ADDRA[10], _4I4426_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_985_9 (_4I4426_$1I4488_$1I4621_ADDRA[9], _4I4426_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_985_8 (_4I4426_$1I4488_$1I4621_ADDRA[8], _4I4426_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_985_7 (_4I4426_$1I4488_$1I4621_ADDRA[7], _4I4426_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_985_6 (_4I4426_$1I4488_$1I4621_ADDRA[6], _4I4426_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_985_5 (_4I4426_$1I4488_$1I4621_ADDRA[5], _4I4426_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_985_4 (_4I4426_$1I4488_$1I4621_ADDRA[4], _4I4426_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_985_3 (_4I4426_$1I4488_$1I4621_ADDRA[3], _4I4426_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_985_2 (_4I4426_$1I4488_$1I4621_ADDRA[2], _4I4426_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_985_1 (_4I4426_$1I4488_$1I4621_ADDRA[1], _4I4426_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_985_0 (_4I4426_$1I4488_$1I4621_ADDRA[0], _4I4426_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _4I4426_$1I4488_$1I4621_ADDRB;
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_986_9 (_4I4426_$1I4488_$1I4621_ADDRB[9], _4I4426_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_986_8 (_4I4426_$1I4488_$1I4621_ADDRB[8], _4I4426_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_986_7 (_4I4426_$1I4488_$1I4621_ADDRB[7], _4I4426_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_986_6 (_4I4426_$1I4488_$1I4621_ADDRB[6], _4I4426_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_986_5 (_4I4426_$1I4488_$1I4621_ADDRB[5], _4I4426_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_986_4 (_4I4426_$1I4488_$1I4621_ADDRB[4], _4I4426_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_986_3 (_4I4426_$1I4488_$1I4621_ADDRB[3], _4I4426_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_986_2 (_4I4426_$1I4488_$1I4621_ADDRB[2], _4I4426_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_986_1 (_4I4426_$1I4488_$1I4621_ADDRB[1], _4I4426_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_986_0 (_4I4426_$1I4488_$1I4621_ADDRB[0], _4I4426_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _4I4426_$1I4488_$1I4621_CLKA;
 reg [1:16] _4I4426_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_987 (_4I4426_$1I4488_$1I4621_CLKA, _4I4426_$1I4488_$1I4621_CLKA__vlIN);

 wire  _4I4426_$1I4488_$1I4621_CLKB;
 reg [1:16] _4I4426_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_988 (_4I4426_$1I4488_$1I4621_CLKB, _4I4426_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _4I4426_$1I4488_$1I4621_DIA;
 reg [1:16] _4I4426_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_989_7 (_4I4426_$1I4488_$1I4621_DIA[7], _4I4426_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_989_6 (_4I4426_$1I4488_$1I4621_DIA[6], _4I4426_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_989_5 (_4I4426_$1I4488_$1I4621_DIA[5], _4I4426_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_989_4 (_4I4426_$1I4488_$1I4621_DIA[4], _4I4426_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_989_3 (_4I4426_$1I4488_$1I4621_DIA[3], _4I4426_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_989_2 (_4I4426_$1I4488_$1I4621_DIA[2], _4I4426_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_989_1 (_4I4426_$1I4488_$1I4621_DIA[1], _4I4426_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_989_0 (_4I4426_$1I4488_$1I4621_DIA[0], _4I4426_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _4I4426_$1I4488_$1I4621_DIB;
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_990_15 (_4I4426_$1I4488_$1I4621_DIB[15], _4I4426_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_990_14 (_4I4426_$1I4488_$1I4621_DIB[14], _4I4426_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_990_13 (_4I4426_$1I4488_$1I4621_DIB[13], _4I4426_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_990_12 (_4I4426_$1I4488_$1I4621_DIB[12], _4I4426_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_990_11 (_4I4426_$1I4488_$1I4621_DIB[11], _4I4426_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_990_10 (_4I4426_$1I4488_$1I4621_DIB[10], _4I4426_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_990_9 (_4I4426_$1I4488_$1I4621_DIB[9], _4I4426_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_990_8 (_4I4426_$1I4488_$1I4621_DIB[8], _4I4426_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_990_7 (_4I4426_$1I4488_$1I4621_DIB[7], _4I4426_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_990_6 (_4I4426_$1I4488_$1I4621_DIB[6], _4I4426_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_990_5 (_4I4426_$1I4488_$1I4621_DIB[5], _4I4426_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_990_4 (_4I4426_$1I4488_$1I4621_DIB[4], _4I4426_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_990_3 (_4I4426_$1I4488_$1I4621_DIB[3], _4I4426_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_990_2 (_4I4426_$1I4488_$1I4621_DIB[2], _4I4426_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_990_1 (_4I4426_$1I4488_$1I4621_DIB[1], _4I4426_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_990_0 (_4I4426_$1I4488_$1I4621_DIB[0], _4I4426_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _4I4426_$1I4488_$1I4621_DIPA;
 reg [1:16] _4I4426_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_991_0 (_4I4426_$1I4488_$1I4621_DIPA[0], _4I4426_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _4I4426_$1I4488_$1I4621_DIPB;
 reg [1:16] _4I4426_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_992_1 (_4I4426_$1I4488_$1I4621_DIPB[1], _4I4426_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_992_0 (_4I4426_$1I4488_$1I4621_DIPB[0], _4I4426_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _4I4426_$1I4488_$1I4621_ENA;
 reg [1:16] _4I4426_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_993 (_4I4426_$1I4488_$1I4621_ENA, _4I4426_$1I4488_$1I4621_ENA__vlIN);

 wire  _4I4426_$1I4488_$1I4621_ENB;
 reg [1:16] _4I4426_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_994 (_4I4426_$1I4488_$1I4621_ENB, _4I4426_$1I4488_$1I4621_ENB__vlIN);

 wire  _4I4426_$1I4488_$1I4621_SSRA;
 reg [1:16] _4I4426_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_995 (_4I4426_$1I4488_$1I4621_SSRA, _4I4426_$1I4488_$1I4621_SSRA__vlIN);

 wire  _4I4426_$1I4488_$1I4621_SSRB;
 reg [1:16] _4I4426_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_996 (_4I4426_$1I4488_$1I4621_SSRB, _4I4426_$1I4488_$1I4621_SSRB__vlIN);

 wire  _4I4426_$1I4488_$1I4621_WEA;
 reg [1:16] _4I4426_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_997 (_4I4426_$1I4488_$1I4621_WEA, _4I4426_$1I4488_$1I4621_WEA__vlIN);

 wire  _4I4426_$1I4488_$1I4621_WEB;
 reg [1:16] _4I4426_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_998 (_4I4426_$1I4488_$1I4621_WEB, _4I4426_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _4I4426_$1I4488_$1I4621 ( _4I4426_$1I4488_$1I4621_DOA , _4I4426_$1I4488_$1I4621_DOB , _4I4426_$1I4488_$1I4621_DOPA , _4I4426_$1I4488_$1I4621_DOPB , _4I4426_$1I4488_$1I4621_ADDRA , _4I4426_$1I4488_$1I4621_ADDRB , _4I4426_$1I4488_$1I4621_CLKA , _4I4426_$1I4488_$1I4621_CLKB , _4I4426_$1I4488_$1I4621_DIA , _4I4426_$1I4488_$1I4621_DIB , _4I4426_$1I4488_$1I4621_DIPA , _4I4426_$1I4488_$1I4621_DIPB , _4I4426_$1I4488_$1I4621_ENA , _4I4426_$1I4488_$1I4621_ENB , _4I4426_$1I4488_$1I4621_SSRA , _4I4426_$1I4488_$1I4621_SSRB , _4I4426_$1I4488_$1I4621_WEA , _4I4426_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4426_$1I4488_$1I4620_DOA;

 wire [15:0] _4I4426_$1I4488_$1I4620_DOB;

 wire [0:0] _4I4426_$1I4488_$1I4620_DOPA;

 wire [1:0] _4I4426_$1I4488_$1I4620_DOPB;

 wire [10:0] _4I4426_$1I4488_$1I4620_ADDRA;
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_999_10 (_4I4426_$1I4488_$1I4620_ADDRA[10], _4I4426_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_999_9 (_4I4426_$1I4488_$1I4620_ADDRA[9], _4I4426_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_999_8 (_4I4426_$1I4488_$1I4620_ADDRA[8], _4I4426_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_999_7 (_4I4426_$1I4488_$1I4620_ADDRA[7], _4I4426_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_999_6 (_4I4426_$1I4488_$1I4620_ADDRA[6], _4I4426_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_999_5 (_4I4426_$1I4488_$1I4620_ADDRA[5], _4I4426_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_999_4 (_4I4426_$1I4488_$1I4620_ADDRA[4], _4I4426_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_999_3 (_4I4426_$1I4488_$1I4620_ADDRA[3], _4I4426_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_999_2 (_4I4426_$1I4488_$1I4620_ADDRA[2], _4I4426_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_999_1 (_4I4426_$1I4488_$1I4620_ADDRA[1], _4I4426_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_999_0 (_4I4426_$1I4488_$1I4620_ADDRA[0], _4I4426_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _4I4426_$1I4488_$1I4620_ADDRB;
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1000_9 (_4I4426_$1I4488_$1I4620_ADDRB[9], _4I4426_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1000_8 (_4I4426_$1I4488_$1I4620_ADDRB[8], _4I4426_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1000_7 (_4I4426_$1I4488_$1I4620_ADDRB[7], _4I4426_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1000_6 (_4I4426_$1I4488_$1I4620_ADDRB[6], _4I4426_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1000_5 (_4I4426_$1I4488_$1I4620_ADDRB[5], _4I4426_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1000_4 (_4I4426_$1I4488_$1I4620_ADDRB[4], _4I4426_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1000_3 (_4I4426_$1I4488_$1I4620_ADDRB[3], _4I4426_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1000_2 (_4I4426_$1I4488_$1I4620_ADDRB[2], _4I4426_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1000_1 (_4I4426_$1I4488_$1I4620_ADDRB[1], _4I4426_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1000_0 (_4I4426_$1I4488_$1I4620_ADDRB[0], _4I4426_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _4I4426_$1I4488_$1I4620_CLKA;
 reg [1:16] _4I4426_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1001 (_4I4426_$1I4488_$1I4620_CLKA, _4I4426_$1I4488_$1I4620_CLKA__vlIN);

 wire  _4I4426_$1I4488_$1I4620_CLKB;
 reg [1:16] _4I4426_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1002 (_4I4426_$1I4488_$1I4620_CLKB, _4I4426_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _4I4426_$1I4488_$1I4620_DIA;
 reg [1:16] _4I4426_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1003_7 (_4I4426_$1I4488_$1I4620_DIA[7], _4I4426_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1003_6 (_4I4426_$1I4488_$1I4620_DIA[6], _4I4426_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1003_5 (_4I4426_$1I4488_$1I4620_DIA[5], _4I4426_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1003_4 (_4I4426_$1I4488_$1I4620_DIA[4], _4I4426_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1003_3 (_4I4426_$1I4488_$1I4620_DIA[3], _4I4426_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1003_2 (_4I4426_$1I4488_$1I4620_DIA[2], _4I4426_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1003_1 (_4I4426_$1I4488_$1I4620_DIA[1], _4I4426_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1003_0 (_4I4426_$1I4488_$1I4620_DIA[0], _4I4426_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _4I4426_$1I4488_$1I4620_DIB;
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1004_15 (_4I4426_$1I4488_$1I4620_DIB[15], _4I4426_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1004_14 (_4I4426_$1I4488_$1I4620_DIB[14], _4I4426_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1004_13 (_4I4426_$1I4488_$1I4620_DIB[13], _4I4426_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1004_12 (_4I4426_$1I4488_$1I4620_DIB[12], _4I4426_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1004_11 (_4I4426_$1I4488_$1I4620_DIB[11], _4I4426_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1004_10 (_4I4426_$1I4488_$1I4620_DIB[10], _4I4426_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1004_9 (_4I4426_$1I4488_$1I4620_DIB[9], _4I4426_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1004_8 (_4I4426_$1I4488_$1I4620_DIB[8], _4I4426_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1004_7 (_4I4426_$1I4488_$1I4620_DIB[7], _4I4426_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1004_6 (_4I4426_$1I4488_$1I4620_DIB[6], _4I4426_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1004_5 (_4I4426_$1I4488_$1I4620_DIB[5], _4I4426_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1004_4 (_4I4426_$1I4488_$1I4620_DIB[4], _4I4426_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1004_3 (_4I4426_$1I4488_$1I4620_DIB[3], _4I4426_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1004_2 (_4I4426_$1I4488_$1I4620_DIB[2], _4I4426_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1004_1 (_4I4426_$1I4488_$1I4620_DIB[1], _4I4426_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1004_0 (_4I4426_$1I4488_$1I4620_DIB[0], _4I4426_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _4I4426_$1I4488_$1I4620_DIPA;
 reg [1:16] _4I4426_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1005_0 (_4I4426_$1I4488_$1I4620_DIPA[0], _4I4426_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _4I4426_$1I4488_$1I4620_DIPB;
 reg [1:16] _4I4426_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1006_1 (_4I4426_$1I4488_$1I4620_DIPB[1], _4I4426_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _4I4426_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1006_0 (_4I4426_$1I4488_$1I4620_DIPB[0], _4I4426_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _4I4426_$1I4488_$1I4620_ENA;
 reg [1:16] _4I4426_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1007 (_4I4426_$1I4488_$1I4620_ENA, _4I4426_$1I4488_$1I4620_ENA__vlIN);

 wire  _4I4426_$1I4488_$1I4620_ENB;
 reg [1:16] _4I4426_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1008 (_4I4426_$1I4488_$1I4620_ENB, _4I4426_$1I4488_$1I4620_ENB__vlIN);

 wire  _4I4426_$1I4488_$1I4620_SSRA;
 reg [1:16] _4I4426_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1009 (_4I4426_$1I4488_$1I4620_SSRA, _4I4426_$1I4488_$1I4620_SSRA__vlIN);

 wire  _4I4426_$1I4488_$1I4620_SSRB;
 reg [1:16] _4I4426_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1010 (_4I4426_$1I4488_$1I4620_SSRB, _4I4426_$1I4488_$1I4620_SSRB__vlIN);

 wire  _4I4426_$1I4488_$1I4620_WEA;
 reg [1:16] _4I4426_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1011 (_4I4426_$1I4488_$1I4620_WEA, _4I4426_$1I4488_$1I4620_WEA__vlIN);

 wire  _4I4426_$1I4488_$1I4620_WEB;
 reg [1:16] _4I4426_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1012 (_4I4426_$1I4488_$1I4620_WEB, _4I4426_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _4I4426_$1I4488_$1I4620 ( _4I4426_$1I4488_$1I4620_DOA , _4I4426_$1I4488_$1I4620_DOB , _4I4426_$1I4488_$1I4620_DOPA , _4I4426_$1I4488_$1I4620_DOPB , _4I4426_$1I4488_$1I4620_ADDRA , _4I4426_$1I4488_$1I4620_ADDRB , _4I4426_$1I4488_$1I4620_CLKA , _4I4426_$1I4488_$1I4620_CLKB , _4I4426_$1I4488_$1I4620_DIA , _4I4426_$1I4488_$1I4620_DIB , _4I4426_$1I4488_$1I4620_DIPA , _4I4426_$1I4488_$1I4620_DIPB , _4I4426_$1I4488_$1I4620_ENA , _4I4426_$1I4488_$1I4620_ENB , _4I4426_$1I4488_$1I4620_SSRA , _4I4426_$1I4488_$1I4620_SSRB , _4I4426_$1I4488_$1I4620_WEA , _4I4426_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4399_$1I4488_$1I4621_DOA;

 wire [15:0] _4I4399_$1I4488_$1I4621_DOB;

 wire [0:0] _4I4399_$1I4488_$1I4621_DOPA;

 wire [1:0] _4I4399_$1I4488_$1I4621_DOPB;

 wire [10:0] _4I4399_$1I4488_$1I4621_ADDRA;
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1013_10 (_4I4399_$1I4488_$1I4621_ADDRA[10], _4I4399_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1013_9 (_4I4399_$1I4488_$1I4621_ADDRA[9], _4I4399_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1013_8 (_4I4399_$1I4488_$1I4621_ADDRA[8], _4I4399_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1013_7 (_4I4399_$1I4488_$1I4621_ADDRA[7], _4I4399_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1013_6 (_4I4399_$1I4488_$1I4621_ADDRA[6], _4I4399_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1013_5 (_4I4399_$1I4488_$1I4621_ADDRA[5], _4I4399_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1013_4 (_4I4399_$1I4488_$1I4621_ADDRA[4], _4I4399_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1013_3 (_4I4399_$1I4488_$1I4621_ADDRA[3], _4I4399_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1013_2 (_4I4399_$1I4488_$1I4621_ADDRA[2], _4I4399_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1013_1 (_4I4399_$1I4488_$1I4621_ADDRA[1], _4I4399_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1013_0 (_4I4399_$1I4488_$1I4621_ADDRA[0], _4I4399_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _4I4399_$1I4488_$1I4621_ADDRB;
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_1014_9 (_4I4399_$1I4488_$1I4621_ADDRB[9], _4I4399_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_1014_8 (_4I4399_$1I4488_$1I4621_ADDRB[8], _4I4399_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_1014_7 (_4I4399_$1I4488_$1I4621_ADDRB[7], _4I4399_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_1014_6 (_4I4399_$1I4488_$1I4621_ADDRB[6], _4I4399_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_1014_5 (_4I4399_$1I4488_$1I4621_ADDRB[5], _4I4399_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_1014_4 (_4I4399_$1I4488_$1I4621_ADDRB[4], _4I4399_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_1014_3 (_4I4399_$1I4488_$1I4621_ADDRB[3], _4I4399_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_1014_2 (_4I4399_$1I4488_$1I4621_ADDRB[2], _4I4399_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_1014_1 (_4I4399_$1I4488_$1I4621_ADDRB[1], _4I4399_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_1014_0 (_4I4399_$1I4488_$1I4621_ADDRB[0], _4I4399_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _4I4399_$1I4488_$1I4621_CLKA;
 reg [1:16] _4I4399_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_1015 (_4I4399_$1I4488_$1I4621_CLKA, _4I4399_$1I4488_$1I4621_CLKA__vlIN);

 wire  _4I4399_$1I4488_$1I4621_CLKB;
 reg [1:16] _4I4399_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_1016 (_4I4399_$1I4488_$1I4621_CLKB, _4I4399_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _4I4399_$1I4488_$1I4621_DIA;
 reg [1:16] _4I4399_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_1017_7 (_4I4399_$1I4488_$1I4621_DIA[7], _4I4399_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_1017_6 (_4I4399_$1I4488_$1I4621_DIA[6], _4I4399_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_1017_5 (_4I4399_$1I4488_$1I4621_DIA[5], _4I4399_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_1017_4 (_4I4399_$1I4488_$1I4621_DIA[4], _4I4399_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_1017_3 (_4I4399_$1I4488_$1I4621_DIA[3], _4I4399_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_1017_2 (_4I4399_$1I4488_$1I4621_DIA[2], _4I4399_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_1017_1 (_4I4399_$1I4488_$1I4621_DIA[1], _4I4399_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_1017_0 (_4I4399_$1I4488_$1I4621_DIA[0], _4I4399_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _4I4399_$1I4488_$1I4621_DIB;
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_1018_15 (_4I4399_$1I4488_$1I4621_DIB[15], _4I4399_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_1018_14 (_4I4399_$1I4488_$1I4621_DIB[14], _4I4399_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_1018_13 (_4I4399_$1I4488_$1I4621_DIB[13], _4I4399_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_1018_12 (_4I4399_$1I4488_$1I4621_DIB[12], _4I4399_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_1018_11 (_4I4399_$1I4488_$1I4621_DIB[11], _4I4399_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_1018_10 (_4I4399_$1I4488_$1I4621_DIB[10], _4I4399_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_1018_9 (_4I4399_$1I4488_$1I4621_DIB[9], _4I4399_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_1018_8 (_4I4399_$1I4488_$1I4621_DIB[8], _4I4399_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_1018_7 (_4I4399_$1I4488_$1I4621_DIB[7], _4I4399_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_1018_6 (_4I4399_$1I4488_$1I4621_DIB[6], _4I4399_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_1018_5 (_4I4399_$1I4488_$1I4621_DIB[5], _4I4399_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_1018_4 (_4I4399_$1I4488_$1I4621_DIB[4], _4I4399_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_1018_3 (_4I4399_$1I4488_$1I4621_DIB[3], _4I4399_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_1018_2 (_4I4399_$1I4488_$1I4621_DIB[2], _4I4399_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_1018_1 (_4I4399_$1I4488_$1I4621_DIB[1], _4I4399_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_1018_0 (_4I4399_$1I4488_$1I4621_DIB[0], _4I4399_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _4I4399_$1I4488_$1I4621_DIPA;
 reg [1:16] _4I4399_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_1019_0 (_4I4399_$1I4488_$1I4621_DIPA[0], _4I4399_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _4I4399_$1I4488_$1I4621_DIPB;
 reg [1:16] _4I4399_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_1020_1 (_4I4399_$1I4488_$1I4621_DIPB[1], _4I4399_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_1020_0 (_4I4399_$1I4488_$1I4621_DIPB[0], _4I4399_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _4I4399_$1I4488_$1I4621_ENA;
 reg [1:16] _4I4399_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_1021 (_4I4399_$1I4488_$1I4621_ENA, _4I4399_$1I4488_$1I4621_ENA__vlIN);

 wire  _4I4399_$1I4488_$1I4621_ENB;
 reg [1:16] _4I4399_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_1022 (_4I4399_$1I4488_$1I4621_ENB, _4I4399_$1I4488_$1I4621_ENB__vlIN);

 wire  _4I4399_$1I4488_$1I4621_SSRA;
 reg [1:16] _4I4399_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_1023 (_4I4399_$1I4488_$1I4621_SSRA, _4I4399_$1I4488_$1I4621_SSRA__vlIN);

 wire  _4I4399_$1I4488_$1I4621_SSRB;
 reg [1:16] _4I4399_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_1024 (_4I4399_$1I4488_$1I4621_SSRB, _4I4399_$1I4488_$1I4621_SSRB__vlIN);

 wire  _4I4399_$1I4488_$1I4621_WEA;
 reg [1:16] _4I4399_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_1025 (_4I4399_$1I4488_$1I4621_WEA, _4I4399_$1I4488_$1I4621_WEA__vlIN);

 wire  _4I4399_$1I4488_$1I4621_WEB;
 reg [1:16] _4I4399_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_1026 (_4I4399_$1I4488_$1I4621_WEB, _4I4399_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _4I4399_$1I4488_$1I4621 ( _4I4399_$1I4488_$1I4621_DOA , _4I4399_$1I4488_$1I4621_DOB , _4I4399_$1I4488_$1I4621_DOPA , _4I4399_$1I4488_$1I4621_DOPB , _4I4399_$1I4488_$1I4621_ADDRA , _4I4399_$1I4488_$1I4621_ADDRB , _4I4399_$1I4488_$1I4621_CLKA , _4I4399_$1I4488_$1I4621_CLKB , _4I4399_$1I4488_$1I4621_DIA , _4I4399_$1I4488_$1I4621_DIB , _4I4399_$1I4488_$1I4621_DIPA , _4I4399_$1I4488_$1I4621_DIPB , _4I4399_$1I4488_$1I4621_ENA , _4I4399_$1I4488_$1I4621_ENB , _4I4399_$1I4488_$1I4621_SSRA , _4I4399_$1I4488_$1I4621_SSRB , _4I4399_$1I4488_$1I4621_WEA , _4I4399_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4399_$1I4488_$1I4620_DOA;

 wire [15:0] _4I4399_$1I4488_$1I4620_DOB;

 wire [0:0] _4I4399_$1I4488_$1I4620_DOPA;

 wire [1:0] _4I4399_$1I4488_$1I4620_DOPB;

 wire [10:0] _4I4399_$1I4488_$1I4620_ADDRA;
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_1027_10 (_4I4399_$1I4488_$1I4620_ADDRA[10], _4I4399_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_1027_9 (_4I4399_$1I4488_$1I4620_ADDRA[9], _4I4399_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_1027_8 (_4I4399_$1I4488_$1I4620_ADDRA[8], _4I4399_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_1027_7 (_4I4399_$1I4488_$1I4620_ADDRA[7], _4I4399_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_1027_6 (_4I4399_$1I4488_$1I4620_ADDRA[6], _4I4399_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_1027_5 (_4I4399_$1I4488_$1I4620_ADDRA[5], _4I4399_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_1027_4 (_4I4399_$1I4488_$1I4620_ADDRA[4], _4I4399_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_1027_3 (_4I4399_$1I4488_$1I4620_ADDRA[3], _4I4399_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_1027_2 (_4I4399_$1I4488_$1I4620_ADDRA[2], _4I4399_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_1027_1 (_4I4399_$1I4488_$1I4620_ADDRA[1], _4I4399_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_1027_0 (_4I4399_$1I4488_$1I4620_ADDRA[0], _4I4399_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _4I4399_$1I4488_$1I4620_ADDRB;
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1028_9 (_4I4399_$1I4488_$1I4620_ADDRB[9], _4I4399_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1028_8 (_4I4399_$1I4488_$1I4620_ADDRB[8], _4I4399_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1028_7 (_4I4399_$1I4488_$1I4620_ADDRB[7], _4I4399_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1028_6 (_4I4399_$1I4488_$1I4620_ADDRB[6], _4I4399_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1028_5 (_4I4399_$1I4488_$1I4620_ADDRB[5], _4I4399_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1028_4 (_4I4399_$1I4488_$1I4620_ADDRB[4], _4I4399_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1028_3 (_4I4399_$1I4488_$1I4620_ADDRB[3], _4I4399_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1028_2 (_4I4399_$1I4488_$1I4620_ADDRB[2], _4I4399_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1028_1 (_4I4399_$1I4488_$1I4620_ADDRB[1], _4I4399_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1028_0 (_4I4399_$1I4488_$1I4620_ADDRB[0], _4I4399_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _4I4399_$1I4488_$1I4620_CLKA;
 reg [1:16] _4I4399_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1029 (_4I4399_$1I4488_$1I4620_CLKA, _4I4399_$1I4488_$1I4620_CLKA__vlIN);

 wire  _4I4399_$1I4488_$1I4620_CLKB;
 reg [1:16] _4I4399_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1030 (_4I4399_$1I4488_$1I4620_CLKB, _4I4399_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _4I4399_$1I4488_$1I4620_DIA;
 reg [1:16] _4I4399_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1031_7 (_4I4399_$1I4488_$1I4620_DIA[7], _4I4399_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1031_6 (_4I4399_$1I4488_$1I4620_DIA[6], _4I4399_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1031_5 (_4I4399_$1I4488_$1I4620_DIA[5], _4I4399_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1031_4 (_4I4399_$1I4488_$1I4620_DIA[4], _4I4399_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1031_3 (_4I4399_$1I4488_$1I4620_DIA[3], _4I4399_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1031_2 (_4I4399_$1I4488_$1I4620_DIA[2], _4I4399_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1031_1 (_4I4399_$1I4488_$1I4620_DIA[1], _4I4399_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1031_0 (_4I4399_$1I4488_$1I4620_DIA[0], _4I4399_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _4I4399_$1I4488_$1I4620_DIB;
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1032_15 (_4I4399_$1I4488_$1I4620_DIB[15], _4I4399_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1032_14 (_4I4399_$1I4488_$1I4620_DIB[14], _4I4399_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1032_13 (_4I4399_$1I4488_$1I4620_DIB[13], _4I4399_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1032_12 (_4I4399_$1I4488_$1I4620_DIB[12], _4I4399_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1032_11 (_4I4399_$1I4488_$1I4620_DIB[11], _4I4399_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1032_10 (_4I4399_$1I4488_$1I4620_DIB[10], _4I4399_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1032_9 (_4I4399_$1I4488_$1I4620_DIB[9], _4I4399_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1032_8 (_4I4399_$1I4488_$1I4620_DIB[8], _4I4399_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1032_7 (_4I4399_$1I4488_$1I4620_DIB[7], _4I4399_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1032_6 (_4I4399_$1I4488_$1I4620_DIB[6], _4I4399_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1032_5 (_4I4399_$1I4488_$1I4620_DIB[5], _4I4399_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1032_4 (_4I4399_$1I4488_$1I4620_DIB[4], _4I4399_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1032_3 (_4I4399_$1I4488_$1I4620_DIB[3], _4I4399_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1032_2 (_4I4399_$1I4488_$1I4620_DIB[2], _4I4399_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1032_1 (_4I4399_$1I4488_$1I4620_DIB[1], _4I4399_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1032_0 (_4I4399_$1I4488_$1I4620_DIB[0], _4I4399_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _4I4399_$1I4488_$1I4620_DIPA;
 reg [1:16] _4I4399_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1033_0 (_4I4399_$1I4488_$1I4620_DIPA[0], _4I4399_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _4I4399_$1I4488_$1I4620_DIPB;
 reg [1:16] _4I4399_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1034_1 (_4I4399_$1I4488_$1I4620_DIPB[1], _4I4399_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _4I4399_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1034_0 (_4I4399_$1I4488_$1I4620_DIPB[0], _4I4399_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _4I4399_$1I4488_$1I4620_ENA;
 reg [1:16] _4I4399_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1035 (_4I4399_$1I4488_$1I4620_ENA, _4I4399_$1I4488_$1I4620_ENA__vlIN);

 wire  _4I4399_$1I4488_$1I4620_ENB;
 reg [1:16] _4I4399_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1036 (_4I4399_$1I4488_$1I4620_ENB, _4I4399_$1I4488_$1I4620_ENB__vlIN);

 wire  _4I4399_$1I4488_$1I4620_SSRA;
 reg [1:16] _4I4399_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1037 (_4I4399_$1I4488_$1I4620_SSRA, _4I4399_$1I4488_$1I4620_SSRA__vlIN);

 wire  _4I4399_$1I4488_$1I4620_SSRB;
 reg [1:16] _4I4399_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1038 (_4I4399_$1I4488_$1I4620_SSRB, _4I4399_$1I4488_$1I4620_SSRB__vlIN);

 wire  _4I4399_$1I4488_$1I4620_WEA;
 reg [1:16] _4I4399_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1039 (_4I4399_$1I4488_$1I4620_WEA, _4I4399_$1I4488_$1I4620_WEA__vlIN);

 wire  _4I4399_$1I4488_$1I4620_WEB;
 reg [1:16] _4I4399_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1040 (_4I4399_$1I4488_$1I4620_WEB, _4I4399_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _4I4399_$1I4488_$1I4620 ( _4I4399_$1I4488_$1I4620_DOA , _4I4399_$1I4488_$1I4620_DOB , _4I4399_$1I4488_$1I4620_DOPA , _4I4399_$1I4488_$1I4620_DOPB , _4I4399_$1I4488_$1I4620_ADDRA , _4I4399_$1I4488_$1I4620_ADDRB , _4I4399_$1I4488_$1I4620_CLKA , _4I4399_$1I4488_$1I4620_CLKB , _4I4399_$1I4488_$1I4620_DIA , _4I4399_$1I4488_$1I4620_DIB , _4I4399_$1I4488_$1I4620_DIPA , _4I4399_$1I4488_$1I4620_DIPB , _4I4399_$1I4488_$1I4620_ENA , _4I4399_$1I4488_$1I4620_ENB , _4I4399_$1I4488_$1I4620_SSRA , _4I4399_$1I4488_$1I4620_SSRB , _4I4399_$1I4488_$1I4620_WEA , _4I4399_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4365_$1I4488_$1I4621_DOA;

 wire [15:0] _4I4365_$1I4488_$1I4621_DOB;

 wire [0:0] _4I4365_$1I4488_$1I4621_DOPA;

 wire [1:0] _4I4365_$1I4488_$1I4621_DOPB;

 wire [10:0] _4I4365_$1I4488_$1I4621_ADDRA;
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1041_10 (_4I4365_$1I4488_$1I4621_ADDRA[10], _4I4365_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1041_9 (_4I4365_$1I4488_$1I4621_ADDRA[9], _4I4365_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1041_8 (_4I4365_$1I4488_$1I4621_ADDRA[8], _4I4365_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1041_7 (_4I4365_$1I4488_$1I4621_ADDRA[7], _4I4365_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1041_6 (_4I4365_$1I4488_$1I4621_ADDRA[6], _4I4365_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1041_5 (_4I4365_$1I4488_$1I4621_ADDRA[5], _4I4365_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1041_4 (_4I4365_$1I4488_$1I4621_ADDRA[4], _4I4365_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1041_3 (_4I4365_$1I4488_$1I4621_ADDRA[3], _4I4365_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1041_2 (_4I4365_$1I4488_$1I4621_ADDRA[2], _4I4365_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1041_1 (_4I4365_$1I4488_$1I4621_ADDRA[1], _4I4365_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1041_0 (_4I4365_$1I4488_$1I4621_ADDRA[0], _4I4365_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _4I4365_$1I4488_$1I4621_ADDRB;
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_1042_9 (_4I4365_$1I4488_$1I4621_ADDRB[9], _4I4365_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_1042_8 (_4I4365_$1I4488_$1I4621_ADDRB[8], _4I4365_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_1042_7 (_4I4365_$1I4488_$1I4621_ADDRB[7], _4I4365_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_1042_6 (_4I4365_$1I4488_$1I4621_ADDRB[6], _4I4365_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_1042_5 (_4I4365_$1I4488_$1I4621_ADDRB[5], _4I4365_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_1042_4 (_4I4365_$1I4488_$1I4621_ADDRB[4], _4I4365_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_1042_3 (_4I4365_$1I4488_$1I4621_ADDRB[3], _4I4365_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_1042_2 (_4I4365_$1I4488_$1I4621_ADDRB[2], _4I4365_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_1042_1 (_4I4365_$1I4488_$1I4621_ADDRB[1], _4I4365_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_1042_0 (_4I4365_$1I4488_$1I4621_ADDRB[0], _4I4365_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _4I4365_$1I4488_$1I4621_CLKA;
 reg [1:16] _4I4365_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_1043 (_4I4365_$1I4488_$1I4621_CLKA, _4I4365_$1I4488_$1I4621_CLKA__vlIN);

 wire  _4I4365_$1I4488_$1I4621_CLKB;
 reg [1:16] _4I4365_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_1044 (_4I4365_$1I4488_$1I4621_CLKB, _4I4365_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _4I4365_$1I4488_$1I4621_DIA;
 reg [1:16] _4I4365_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_1045_7 (_4I4365_$1I4488_$1I4621_DIA[7], _4I4365_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_1045_6 (_4I4365_$1I4488_$1I4621_DIA[6], _4I4365_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_1045_5 (_4I4365_$1I4488_$1I4621_DIA[5], _4I4365_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_1045_4 (_4I4365_$1I4488_$1I4621_DIA[4], _4I4365_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_1045_3 (_4I4365_$1I4488_$1I4621_DIA[3], _4I4365_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_1045_2 (_4I4365_$1I4488_$1I4621_DIA[2], _4I4365_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_1045_1 (_4I4365_$1I4488_$1I4621_DIA[1], _4I4365_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_1045_0 (_4I4365_$1I4488_$1I4621_DIA[0], _4I4365_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _4I4365_$1I4488_$1I4621_DIB;
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_1046_15 (_4I4365_$1I4488_$1I4621_DIB[15], _4I4365_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_1046_14 (_4I4365_$1I4488_$1I4621_DIB[14], _4I4365_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_1046_13 (_4I4365_$1I4488_$1I4621_DIB[13], _4I4365_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_1046_12 (_4I4365_$1I4488_$1I4621_DIB[12], _4I4365_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_1046_11 (_4I4365_$1I4488_$1I4621_DIB[11], _4I4365_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_1046_10 (_4I4365_$1I4488_$1I4621_DIB[10], _4I4365_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_1046_9 (_4I4365_$1I4488_$1I4621_DIB[9], _4I4365_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_1046_8 (_4I4365_$1I4488_$1I4621_DIB[8], _4I4365_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_1046_7 (_4I4365_$1I4488_$1I4621_DIB[7], _4I4365_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_1046_6 (_4I4365_$1I4488_$1I4621_DIB[6], _4I4365_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_1046_5 (_4I4365_$1I4488_$1I4621_DIB[5], _4I4365_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_1046_4 (_4I4365_$1I4488_$1I4621_DIB[4], _4I4365_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_1046_3 (_4I4365_$1I4488_$1I4621_DIB[3], _4I4365_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_1046_2 (_4I4365_$1I4488_$1I4621_DIB[2], _4I4365_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_1046_1 (_4I4365_$1I4488_$1I4621_DIB[1], _4I4365_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_1046_0 (_4I4365_$1I4488_$1I4621_DIB[0], _4I4365_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _4I4365_$1I4488_$1I4621_DIPA;
 reg [1:16] _4I4365_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_1047_0 (_4I4365_$1I4488_$1I4621_DIPA[0], _4I4365_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _4I4365_$1I4488_$1I4621_DIPB;
 reg [1:16] _4I4365_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_1048_1 (_4I4365_$1I4488_$1I4621_DIPB[1], _4I4365_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_1048_0 (_4I4365_$1I4488_$1I4621_DIPB[0], _4I4365_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _4I4365_$1I4488_$1I4621_ENA;
 reg [1:16] _4I4365_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_1049 (_4I4365_$1I4488_$1I4621_ENA, _4I4365_$1I4488_$1I4621_ENA__vlIN);

 wire  _4I4365_$1I4488_$1I4621_ENB;
 reg [1:16] _4I4365_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_1050 (_4I4365_$1I4488_$1I4621_ENB, _4I4365_$1I4488_$1I4621_ENB__vlIN);

 wire  _4I4365_$1I4488_$1I4621_SSRA;
 reg [1:16] _4I4365_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_1051 (_4I4365_$1I4488_$1I4621_SSRA, _4I4365_$1I4488_$1I4621_SSRA__vlIN);

 wire  _4I4365_$1I4488_$1I4621_SSRB;
 reg [1:16] _4I4365_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_1052 (_4I4365_$1I4488_$1I4621_SSRB, _4I4365_$1I4488_$1I4621_SSRB__vlIN);

 wire  _4I4365_$1I4488_$1I4621_WEA;
 reg [1:16] _4I4365_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_1053 (_4I4365_$1I4488_$1I4621_WEA, _4I4365_$1I4488_$1I4621_WEA__vlIN);

 wire  _4I4365_$1I4488_$1I4621_WEB;
 reg [1:16] _4I4365_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_1054 (_4I4365_$1I4488_$1I4621_WEB, _4I4365_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _4I4365_$1I4488_$1I4621 ( _4I4365_$1I4488_$1I4621_DOA , _4I4365_$1I4488_$1I4621_DOB , _4I4365_$1I4488_$1I4621_DOPA , _4I4365_$1I4488_$1I4621_DOPB , _4I4365_$1I4488_$1I4621_ADDRA , _4I4365_$1I4488_$1I4621_ADDRB , _4I4365_$1I4488_$1I4621_CLKA , _4I4365_$1I4488_$1I4621_CLKB , _4I4365_$1I4488_$1I4621_DIA , _4I4365_$1I4488_$1I4621_DIB , _4I4365_$1I4488_$1I4621_DIPA , _4I4365_$1I4488_$1I4621_DIPB , _4I4365_$1I4488_$1I4621_ENA , _4I4365_$1I4488_$1I4621_ENB , _4I4365_$1I4488_$1I4621_SSRA , _4I4365_$1I4488_$1I4621_SSRB , _4I4365_$1I4488_$1I4621_WEA , _4I4365_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4365_$1I4488_$1I4620_DOA;

 wire [15:0] _4I4365_$1I4488_$1I4620_DOB;

 wire [0:0] _4I4365_$1I4488_$1I4620_DOPA;

 wire [1:0] _4I4365_$1I4488_$1I4620_DOPB;

 wire [10:0] _4I4365_$1I4488_$1I4620_ADDRA;
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_1055_10 (_4I4365_$1I4488_$1I4620_ADDRA[10], _4I4365_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_1055_9 (_4I4365_$1I4488_$1I4620_ADDRA[9], _4I4365_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_1055_8 (_4I4365_$1I4488_$1I4620_ADDRA[8], _4I4365_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_1055_7 (_4I4365_$1I4488_$1I4620_ADDRA[7], _4I4365_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_1055_6 (_4I4365_$1I4488_$1I4620_ADDRA[6], _4I4365_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_1055_5 (_4I4365_$1I4488_$1I4620_ADDRA[5], _4I4365_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_1055_4 (_4I4365_$1I4488_$1I4620_ADDRA[4], _4I4365_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_1055_3 (_4I4365_$1I4488_$1I4620_ADDRA[3], _4I4365_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_1055_2 (_4I4365_$1I4488_$1I4620_ADDRA[2], _4I4365_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_1055_1 (_4I4365_$1I4488_$1I4620_ADDRA[1], _4I4365_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_1055_0 (_4I4365_$1I4488_$1I4620_ADDRA[0], _4I4365_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _4I4365_$1I4488_$1I4620_ADDRB;
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1056_9 (_4I4365_$1I4488_$1I4620_ADDRB[9], _4I4365_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1056_8 (_4I4365_$1I4488_$1I4620_ADDRB[8], _4I4365_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1056_7 (_4I4365_$1I4488_$1I4620_ADDRB[7], _4I4365_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1056_6 (_4I4365_$1I4488_$1I4620_ADDRB[6], _4I4365_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1056_5 (_4I4365_$1I4488_$1I4620_ADDRB[5], _4I4365_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1056_4 (_4I4365_$1I4488_$1I4620_ADDRB[4], _4I4365_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1056_3 (_4I4365_$1I4488_$1I4620_ADDRB[3], _4I4365_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1056_2 (_4I4365_$1I4488_$1I4620_ADDRB[2], _4I4365_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1056_1 (_4I4365_$1I4488_$1I4620_ADDRB[1], _4I4365_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1056_0 (_4I4365_$1I4488_$1I4620_ADDRB[0], _4I4365_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _4I4365_$1I4488_$1I4620_CLKA;
 reg [1:16] _4I4365_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1057 (_4I4365_$1I4488_$1I4620_CLKA, _4I4365_$1I4488_$1I4620_CLKA__vlIN);

 wire  _4I4365_$1I4488_$1I4620_CLKB;
 reg [1:16] _4I4365_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1058 (_4I4365_$1I4488_$1I4620_CLKB, _4I4365_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _4I4365_$1I4488_$1I4620_DIA;
 reg [1:16] _4I4365_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1059_7 (_4I4365_$1I4488_$1I4620_DIA[7], _4I4365_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1059_6 (_4I4365_$1I4488_$1I4620_DIA[6], _4I4365_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1059_5 (_4I4365_$1I4488_$1I4620_DIA[5], _4I4365_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1059_4 (_4I4365_$1I4488_$1I4620_DIA[4], _4I4365_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1059_3 (_4I4365_$1I4488_$1I4620_DIA[3], _4I4365_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1059_2 (_4I4365_$1I4488_$1I4620_DIA[2], _4I4365_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1059_1 (_4I4365_$1I4488_$1I4620_DIA[1], _4I4365_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1059_0 (_4I4365_$1I4488_$1I4620_DIA[0], _4I4365_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _4I4365_$1I4488_$1I4620_DIB;
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1060_15 (_4I4365_$1I4488_$1I4620_DIB[15], _4I4365_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1060_14 (_4I4365_$1I4488_$1I4620_DIB[14], _4I4365_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1060_13 (_4I4365_$1I4488_$1I4620_DIB[13], _4I4365_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1060_12 (_4I4365_$1I4488_$1I4620_DIB[12], _4I4365_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1060_11 (_4I4365_$1I4488_$1I4620_DIB[11], _4I4365_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1060_10 (_4I4365_$1I4488_$1I4620_DIB[10], _4I4365_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1060_9 (_4I4365_$1I4488_$1I4620_DIB[9], _4I4365_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1060_8 (_4I4365_$1I4488_$1I4620_DIB[8], _4I4365_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1060_7 (_4I4365_$1I4488_$1I4620_DIB[7], _4I4365_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1060_6 (_4I4365_$1I4488_$1I4620_DIB[6], _4I4365_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1060_5 (_4I4365_$1I4488_$1I4620_DIB[5], _4I4365_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1060_4 (_4I4365_$1I4488_$1I4620_DIB[4], _4I4365_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1060_3 (_4I4365_$1I4488_$1I4620_DIB[3], _4I4365_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1060_2 (_4I4365_$1I4488_$1I4620_DIB[2], _4I4365_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1060_1 (_4I4365_$1I4488_$1I4620_DIB[1], _4I4365_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1060_0 (_4I4365_$1I4488_$1I4620_DIB[0], _4I4365_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _4I4365_$1I4488_$1I4620_DIPA;
 reg [1:16] _4I4365_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1061_0 (_4I4365_$1I4488_$1I4620_DIPA[0], _4I4365_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _4I4365_$1I4488_$1I4620_DIPB;
 reg [1:16] _4I4365_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1062_1 (_4I4365_$1I4488_$1I4620_DIPB[1], _4I4365_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _4I4365_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1062_0 (_4I4365_$1I4488_$1I4620_DIPB[0], _4I4365_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _4I4365_$1I4488_$1I4620_ENA;
 reg [1:16] _4I4365_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1063 (_4I4365_$1I4488_$1I4620_ENA, _4I4365_$1I4488_$1I4620_ENA__vlIN);

 wire  _4I4365_$1I4488_$1I4620_ENB;
 reg [1:16] _4I4365_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1064 (_4I4365_$1I4488_$1I4620_ENB, _4I4365_$1I4488_$1I4620_ENB__vlIN);

 wire  _4I4365_$1I4488_$1I4620_SSRA;
 reg [1:16] _4I4365_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1065 (_4I4365_$1I4488_$1I4620_SSRA, _4I4365_$1I4488_$1I4620_SSRA__vlIN);

 wire  _4I4365_$1I4488_$1I4620_SSRB;
 reg [1:16] _4I4365_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1066 (_4I4365_$1I4488_$1I4620_SSRB, _4I4365_$1I4488_$1I4620_SSRB__vlIN);

 wire  _4I4365_$1I4488_$1I4620_WEA;
 reg [1:16] _4I4365_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1067 (_4I4365_$1I4488_$1I4620_WEA, _4I4365_$1I4488_$1I4620_WEA__vlIN);

 wire  _4I4365_$1I4488_$1I4620_WEB;
 reg [1:16] _4I4365_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1068 (_4I4365_$1I4488_$1I4620_WEB, _4I4365_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _4I4365_$1I4488_$1I4620 ( _4I4365_$1I4488_$1I4620_DOA , _4I4365_$1I4488_$1I4620_DOB , _4I4365_$1I4488_$1I4620_DOPA , _4I4365_$1I4488_$1I4620_DOPB , _4I4365_$1I4488_$1I4620_ADDRA , _4I4365_$1I4488_$1I4620_ADDRB , _4I4365_$1I4488_$1I4620_CLKA , _4I4365_$1I4488_$1I4620_CLKB , _4I4365_$1I4488_$1I4620_DIA , _4I4365_$1I4488_$1I4620_DIB , _4I4365_$1I4488_$1I4620_DIPA , _4I4365_$1I4488_$1I4620_DIPB , _4I4365_$1I4488_$1I4620_ENA , _4I4365_$1I4488_$1I4620_ENB , _4I4365_$1I4488_$1I4620_SSRA , _4I4365_$1I4488_$1I4620_SSRB , _4I4365_$1I4488_$1I4620_WEA , _4I4365_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4329_$1I4488_$1I4621_DOA;

 wire [15:0] _4I4329_$1I4488_$1I4621_DOB;

 wire [0:0] _4I4329_$1I4488_$1I4621_DOPA;

 wire [1:0] _4I4329_$1I4488_$1I4621_DOPB;

 wire [10:0] _4I4329_$1I4488_$1I4621_ADDRA;
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1069_10 (_4I4329_$1I4488_$1I4621_ADDRA[10], _4I4329_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1069_9 (_4I4329_$1I4488_$1I4621_ADDRA[9], _4I4329_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1069_8 (_4I4329_$1I4488_$1I4621_ADDRA[8], _4I4329_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1069_7 (_4I4329_$1I4488_$1I4621_ADDRA[7], _4I4329_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1069_6 (_4I4329_$1I4488_$1I4621_ADDRA[6], _4I4329_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1069_5 (_4I4329_$1I4488_$1I4621_ADDRA[5], _4I4329_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1069_4 (_4I4329_$1I4488_$1I4621_ADDRA[4], _4I4329_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1069_3 (_4I4329_$1I4488_$1I4621_ADDRA[3], _4I4329_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1069_2 (_4I4329_$1I4488_$1I4621_ADDRA[2], _4I4329_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1069_1 (_4I4329_$1I4488_$1I4621_ADDRA[1], _4I4329_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1069_0 (_4I4329_$1I4488_$1I4621_ADDRA[0], _4I4329_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _4I4329_$1I4488_$1I4621_ADDRB;
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_1070_9 (_4I4329_$1I4488_$1I4621_ADDRB[9], _4I4329_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_1070_8 (_4I4329_$1I4488_$1I4621_ADDRB[8], _4I4329_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_1070_7 (_4I4329_$1I4488_$1I4621_ADDRB[7], _4I4329_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_1070_6 (_4I4329_$1I4488_$1I4621_ADDRB[6], _4I4329_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_1070_5 (_4I4329_$1I4488_$1I4621_ADDRB[5], _4I4329_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_1070_4 (_4I4329_$1I4488_$1I4621_ADDRB[4], _4I4329_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_1070_3 (_4I4329_$1I4488_$1I4621_ADDRB[3], _4I4329_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_1070_2 (_4I4329_$1I4488_$1I4621_ADDRB[2], _4I4329_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_1070_1 (_4I4329_$1I4488_$1I4621_ADDRB[1], _4I4329_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_1070_0 (_4I4329_$1I4488_$1I4621_ADDRB[0], _4I4329_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _4I4329_$1I4488_$1I4621_CLKA;
 reg [1:16] _4I4329_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_1071 (_4I4329_$1I4488_$1I4621_CLKA, _4I4329_$1I4488_$1I4621_CLKA__vlIN);

 wire  _4I4329_$1I4488_$1I4621_CLKB;
 reg [1:16] _4I4329_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_1072 (_4I4329_$1I4488_$1I4621_CLKB, _4I4329_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _4I4329_$1I4488_$1I4621_DIA;
 reg [1:16] _4I4329_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_1073_7 (_4I4329_$1I4488_$1I4621_DIA[7], _4I4329_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_1073_6 (_4I4329_$1I4488_$1I4621_DIA[6], _4I4329_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_1073_5 (_4I4329_$1I4488_$1I4621_DIA[5], _4I4329_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_1073_4 (_4I4329_$1I4488_$1I4621_DIA[4], _4I4329_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_1073_3 (_4I4329_$1I4488_$1I4621_DIA[3], _4I4329_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_1073_2 (_4I4329_$1I4488_$1I4621_DIA[2], _4I4329_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_1073_1 (_4I4329_$1I4488_$1I4621_DIA[1], _4I4329_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_1073_0 (_4I4329_$1I4488_$1I4621_DIA[0], _4I4329_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _4I4329_$1I4488_$1I4621_DIB;
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_1074_15 (_4I4329_$1I4488_$1I4621_DIB[15], _4I4329_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_1074_14 (_4I4329_$1I4488_$1I4621_DIB[14], _4I4329_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_1074_13 (_4I4329_$1I4488_$1I4621_DIB[13], _4I4329_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_1074_12 (_4I4329_$1I4488_$1I4621_DIB[12], _4I4329_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_1074_11 (_4I4329_$1I4488_$1I4621_DIB[11], _4I4329_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_1074_10 (_4I4329_$1I4488_$1I4621_DIB[10], _4I4329_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_1074_9 (_4I4329_$1I4488_$1I4621_DIB[9], _4I4329_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_1074_8 (_4I4329_$1I4488_$1I4621_DIB[8], _4I4329_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_1074_7 (_4I4329_$1I4488_$1I4621_DIB[7], _4I4329_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_1074_6 (_4I4329_$1I4488_$1I4621_DIB[6], _4I4329_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_1074_5 (_4I4329_$1I4488_$1I4621_DIB[5], _4I4329_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_1074_4 (_4I4329_$1I4488_$1I4621_DIB[4], _4I4329_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_1074_3 (_4I4329_$1I4488_$1I4621_DIB[3], _4I4329_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_1074_2 (_4I4329_$1I4488_$1I4621_DIB[2], _4I4329_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_1074_1 (_4I4329_$1I4488_$1I4621_DIB[1], _4I4329_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_1074_0 (_4I4329_$1I4488_$1I4621_DIB[0], _4I4329_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _4I4329_$1I4488_$1I4621_DIPA;
 reg [1:16] _4I4329_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_1075_0 (_4I4329_$1I4488_$1I4621_DIPA[0], _4I4329_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _4I4329_$1I4488_$1I4621_DIPB;
 reg [1:16] _4I4329_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_1076_1 (_4I4329_$1I4488_$1I4621_DIPB[1], _4I4329_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_1076_0 (_4I4329_$1I4488_$1I4621_DIPB[0], _4I4329_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _4I4329_$1I4488_$1I4621_ENA;
 reg [1:16] _4I4329_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_1077 (_4I4329_$1I4488_$1I4621_ENA, _4I4329_$1I4488_$1I4621_ENA__vlIN);

 wire  _4I4329_$1I4488_$1I4621_ENB;
 reg [1:16] _4I4329_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_1078 (_4I4329_$1I4488_$1I4621_ENB, _4I4329_$1I4488_$1I4621_ENB__vlIN);

 wire  _4I4329_$1I4488_$1I4621_SSRA;
 reg [1:16] _4I4329_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_1079 (_4I4329_$1I4488_$1I4621_SSRA, _4I4329_$1I4488_$1I4621_SSRA__vlIN);

 wire  _4I4329_$1I4488_$1I4621_SSRB;
 reg [1:16] _4I4329_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_1080 (_4I4329_$1I4488_$1I4621_SSRB, _4I4329_$1I4488_$1I4621_SSRB__vlIN);

 wire  _4I4329_$1I4488_$1I4621_WEA;
 reg [1:16] _4I4329_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_1081 (_4I4329_$1I4488_$1I4621_WEA, _4I4329_$1I4488_$1I4621_WEA__vlIN);

 wire  _4I4329_$1I4488_$1I4621_WEB;
 reg [1:16] _4I4329_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_1082 (_4I4329_$1I4488_$1I4621_WEB, _4I4329_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _4I4329_$1I4488_$1I4621 ( _4I4329_$1I4488_$1I4621_DOA , _4I4329_$1I4488_$1I4621_DOB , _4I4329_$1I4488_$1I4621_DOPA , _4I4329_$1I4488_$1I4621_DOPB , _4I4329_$1I4488_$1I4621_ADDRA , _4I4329_$1I4488_$1I4621_ADDRB , _4I4329_$1I4488_$1I4621_CLKA , _4I4329_$1I4488_$1I4621_CLKB , _4I4329_$1I4488_$1I4621_DIA , _4I4329_$1I4488_$1I4621_DIB , _4I4329_$1I4488_$1I4621_DIPA , _4I4329_$1I4488_$1I4621_DIPB , _4I4329_$1I4488_$1I4621_ENA , _4I4329_$1I4488_$1I4621_ENB , _4I4329_$1I4488_$1I4621_SSRA , _4I4329_$1I4488_$1I4621_SSRB , _4I4329_$1I4488_$1I4621_WEA , _4I4329_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _4I4329_$1I4488_$1I4620_DOA;

 wire [15:0] _4I4329_$1I4488_$1I4620_DOB;

 wire [0:0] _4I4329_$1I4488_$1I4620_DOPA;

 wire [1:0] _4I4329_$1I4488_$1I4620_DOPB;

 wire [10:0] _4I4329_$1I4488_$1I4620_ADDRA;
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_1083_10 (_4I4329_$1I4488_$1I4620_ADDRA[10], _4I4329_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_1083_9 (_4I4329_$1I4488_$1I4620_ADDRA[9], _4I4329_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_1083_8 (_4I4329_$1I4488_$1I4620_ADDRA[8], _4I4329_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_1083_7 (_4I4329_$1I4488_$1I4620_ADDRA[7], _4I4329_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_1083_6 (_4I4329_$1I4488_$1I4620_ADDRA[6], _4I4329_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_1083_5 (_4I4329_$1I4488_$1I4620_ADDRA[5], _4I4329_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_1083_4 (_4I4329_$1I4488_$1I4620_ADDRA[4], _4I4329_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_1083_3 (_4I4329_$1I4488_$1I4620_ADDRA[3], _4I4329_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_1083_2 (_4I4329_$1I4488_$1I4620_ADDRA[2], _4I4329_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_1083_1 (_4I4329_$1I4488_$1I4620_ADDRA[1], _4I4329_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_1083_0 (_4I4329_$1I4488_$1I4620_ADDRA[0], _4I4329_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _4I4329_$1I4488_$1I4620_ADDRB;
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1084_9 (_4I4329_$1I4488_$1I4620_ADDRB[9], _4I4329_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1084_8 (_4I4329_$1I4488_$1I4620_ADDRB[8], _4I4329_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1084_7 (_4I4329_$1I4488_$1I4620_ADDRB[7], _4I4329_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1084_6 (_4I4329_$1I4488_$1I4620_ADDRB[6], _4I4329_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1084_5 (_4I4329_$1I4488_$1I4620_ADDRB[5], _4I4329_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1084_4 (_4I4329_$1I4488_$1I4620_ADDRB[4], _4I4329_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1084_3 (_4I4329_$1I4488_$1I4620_ADDRB[3], _4I4329_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1084_2 (_4I4329_$1I4488_$1I4620_ADDRB[2], _4I4329_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1084_1 (_4I4329_$1I4488_$1I4620_ADDRB[1], _4I4329_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1084_0 (_4I4329_$1I4488_$1I4620_ADDRB[0], _4I4329_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _4I4329_$1I4488_$1I4620_CLKA;
 reg [1:16] _4I4329_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1085 (_4I4329_$1I4488_$1I4620_CLKA, _4I4329_$1I4488_$1I4620_CLKA__vlIN);

 wire  _4I4329_$1I4488_$1I4620_CLKB;
 reg [1:16] _4I4329_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1086 (_4I4329_$1I4488_$1I4620_CLKB, _4I4329_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _4I4329_$1I4488_$1I4620_DIA;
 reg [1:16] _4I4329_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1087_7 (_4I4329_$1I4488_$1I4620_DIA[7], _4I4329_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1087_6 (_4I4329_$1I4488_$1I4620_DIA[6], _4I4329_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1087_5 (_4I4329_$1I4488_$1I4620_DIA[5], _4I4329_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1087_4 (_4I4329_$1I4488_$1I4620_DIA[4], _4I4329_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1087_3 (_4I4329_$1I4488_$1I4620_DIA[3], _4I4329_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1087_2 (_4I4329_$1I4488_$1I4620_DIA[2], _4I4329_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1087_1 (_4I4329_$1I4488_$1I4620_DIA[1], _4I4329_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1087_0 (_4I4329_$1I4488_$1I4620_DIA[0], _4I4329_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _4I4329_$1I4488_$1I4620_DIB;
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1088_15 (_4I4329_$1I4488_$1I4620_DIB[15], _4I4329_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1088_14 (_4I4329_$1I4488_$1I4620_DIB[14], _4I4329_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1088_13 (_4I4329_$1I4488_$1I4620_DIB[13], _4I4329_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1088_12 (_4I4329_$1I4488_$1I4620_DIB[12], _4I4329_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1088_11 (_4I4329_$1I4488_$1I4620_DIB[11], _4I4329_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1088_10 (_4I4329_$1I4488_$1I4620_DIB[10], _4I4329_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1088_9 (_4I4329_$1I4488_$1I4620_DIB[9], _4I4329_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1088_8 (_4I4329_$1I4488_$1I4620_DIB[8], _4I4329_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1088_7 (_4I4329_$1I4488_$1I4620_DIB[7], _4I4329_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1088_6 (_4I4329_$1I4488_$1I4620_DIB[6], _4I4329_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1088_5 (_4I4329_$1I4488_$1I4620_DIB[5], _4I4329_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1088_4 (_4I4329_$1I4488_$1I4620_DIB[4], _4I4329_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1088_3 (_4I4329_$1I4488_$1I4620_DIB[3], _4I4329_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1088_2 (_4I4329_$1I4488_$1I4620_DIB[2], _4I4329_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1088_1 (_4I4329_$1I4488_$1I4620_DIB[1], _4I4329_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1088_0 (_4I4329_$1I4488_$1I4620_DIB[0], _4I4329_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _4I4329_$1I4488_$1I4620_DIPA;
 reg [1:16] _4I4329_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1089_0 (_4I4329_$1I4488_$1I4620_DIPA[0], _4I4329_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _4I4329_$1I4488_$1I4620_DIPB;
 reg [1:16] _4I4329_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1090_1 (_4I4329_$1I4488_$1I4620_DIPB[1], _4I4329_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _4I4329_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1090_0 (_4I4329_$1I4488_$1I4620_DIPB[0], _4I4329_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _4I4329_$1I4488_$1I4620_ENA;
 reg [1:16] _4I4329_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1091 (_4I4329_$1I4488_$1I4620_ENA, _4I4329_$1I4488_$1I4620_ENA__vlIN);

 wire  _4I4329_$1I4488_$1I4620_ENB;
 reg [1:16] _4I4329_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1092 (_4I4329_$1I4488_$1I4620_ENB, _4I4329_$1I4488_$1I4620_ENB__vlIN);

 wire  _4I4329_$1I4488_$1I4620_SSRA;
 reg [1:16] _4I4329_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1093 (_4I4329_$1I4488_$1I4620_SSRA, _4I4329_$1I4488_$1I4620_SSRA__vlIN);

 wire  _4I4329_$1I4488_$1I4620_SSRB;
 reg [1:16] _4I4329_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1094 (_4I4329_$1I4488_$1I4620_SSRB, _4I4329_$1I4488_$1I4620_SSRB__vlIN);

 wire  _4I4329_$1I4488_$1I4620_WEA;
 reg [1:16] _4I4329_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1095 (_4I4329_$1I4488_$1I4620_WEA, _4I4329_$1I4488_$1I4620_WEA__vlIN);

 wire  _4I4329_$1I4488_$1I4620_WEB;
 reg [1:16] _4I4329_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1096 (_4I4329_$1I4488_$1I4620_WEB, _4I4329_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _4I4329_$1I4488_$1I4620 ( _4I4329_$1I4488_$1I4620_DOA , _4I4329_$1I4488_$1I4620_DOB , _4I4329_$1I4488_$1I4620_DOPA , _4I4329_$1I4488_$1I4620_DOPB , _4I4329_$1I4488_$1I4620_ADDRA , _4I4329_$1I4488_$1I4620_ADDRB , _4I4329_$1I4488_$1I4620_CLKA , _4I4329_$1I4488_$1I4620_CLKB , _4I4329_$1I4488_$1I4620_DIA , _4I4329_$1I4488_$1I4620_DIB , _4I4329_$1I4488_$1I4620_DIPA , _4I4329_$1I4488_$1I4620_DIPB , _4I4329_$1I4488_$1I4620_ENA , _4I4329_$1I4488_$1I4620_ENB , _4I4329_$1I4488_$1I4620_SSRA , _4I4329_$1I4488_$1I4620_SSRB , _4I4329_$1I4488_$1I4620_WEA , _4I4329_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4551_$1I4488_$1I4621_DOA;

 wire [15:0] _3I4551_$1I4488_$1I4621_DOB;

 wire [0:0] _3I4551_$1I4488_$1I4621_DOPA;

 wire [1:0] _3I4551_$1I4488_$1I4621_DOPB;

 wire [10:0] _3I4551_$1I4488_$1I4621_ADDRA;
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1097_10 (_3I4551_$1I4488_$1I4621_ADDRA[10], _3I4551_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1097_9 (_3I4551_$1I4488_$1I4621_ADDRA[9], _3I4551_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1097_8 (_3I4551_$1I4488_$1I4621_ADDRA[8], _3I4551_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1097_7 (_3I4551_$1I4488_$1I4621_ADDRA[7], _3I4551_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1097_6 (_3I4551_$1I4488_$1I4621_ADDRA[6], _3I4551_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1097_5 (_3I4551_$1I4488_$1I4621_ADDRA[5], _3I4551_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1097_4 (_3I4551_$1I4488_$1I4621_ADDRA[4], _3I4551_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1097_3 (_3I4551_$1I4488_$1I4621_ADDRA[3], _3I4551_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1097_2 (_3I4551_$1I4488_$1I4621_ADDRA[2], _3I4551_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1097_1 (_3I4551_$1I4488_$1I4621_ADDRA[1], _3I4551_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1097_0 (_3I4551_$1I4488_$1I4621_ADDRA[0], _3I4551_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _3I4551_$1I4488_$1I4621_ADDRB;
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_1098_9 (_3I4551_$1I4488_$1I4621_ADDRB[9], _3I4551_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_1098_8 (_3I4551_$1I4488_$1I4621_ADDRB[8], _3I4551_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_1098_7 (_3I4551_$1I4488_$1I4621_ADDRB[7], _3I4551_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_1098_6 (_3I4551_$1I4488_$1I4621_ADDRB[6], _3I4551_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_1098_5 (_3I4551_$1I4488_$1I4621_ADDRB[5], _3I4551_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_1098_4 (_3I4551_$1I4488_$1I4621_ADDRB[4], _3I4551_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_1098_3 (_3I4551_$1I4488_$1I4621_ADDRB[3], _3I4551_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_1098_2 (_3I4551_$1I4488_$1I4621_ADDRB[2], _3I4551_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_1098_1 (_3I4551_$1I4488_$1I4621_ADDRB[1], _3I4551_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_1098_0 (_3I4551_$1I4488_$1I4621_ADDRB[0], _3I4551_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _3I4551_$1I4488_$1I4621_CLKA;
 reg [1:16] _3I4551_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_1099 (_3I4551_$1I4488_$1I4621_CLKA, _3I4551_$1I4488_$1I4621_CLKA__vlIN);

 wire  _3I4551_$1I4488_$1I4621_CLKB;
 reg [1:16] _3I4551_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_1100 (_3I4551_$1I4488_$1I4621_CLKB, _3I4551_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _3I4551_$1I4488_$1I4621_DIA;
 reg [1:16] _3I4551_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_1101_7 (_3I4551_$1I4488_$1I4621_DIA[7], _3I4551_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_1101_6 (_3I4551_$1I4488_$1I4621_DIA[6], _3I4551_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_1101_5 (_3I4551_$1I4488_$1I4621_DIA[5], _3I4551_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_1101_4 (_3I4551_$1I4488_$1I4621_DIA[4], _3I4551_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_1101_3 (_3I4551_$1I4488_$1I4621_DIA[3], _3I4551_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_1101_2 (_3I4551_$1I4488_$1I4621_DIA[2], _3I4551_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_1101_1 (_3I4551_$1I4488_$1I4621_DIA[1], _3I4551_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_1101_0 (_3I4551_$1I4488_$1I4621_DIA[0], _3I4551_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _3I4551_$1I4488_$1I4621_DIB;
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_1102_15 (_3I4551_$1I4488_$1I4621_DIB[15], _3I4551_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_1102_14 (_3I4551_$1I4488_$1I4621_DIB[14], _3I4551_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_1102_13 (_3I4551_$1I4488_$1I4621_DIB[13], _3I4551_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_1102_12 (_3I4551_$1I4488_$1I4621_DIB[12], _3I4551_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_1102_11 (_3I4551_$1I4488_$1I4621_DIB[11], _3I4551_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_1102_10 (_3I4551_$1I4488_$1I4621_DIB[10], _3I4551_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_1102_9 (_3I4551_$1I4488_$1I4621_DIB[9], _3I4551_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_1102_8 (_3I4551_$1I4488_$1I4621_DIB[8], _3I4551_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_1102_7 (_3I4551_$1I4488_$1I4621_DIB[7], _3I4551_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_1102_6 (_3I4551_$1I4488_$1I4621_DIB[6], _3I4551_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_1102_5 (_3I4551_$1I4488_$1I4621_DIB[5], _3I4551_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_1102_4 (_3I4551_$1I4488_$1I4621_DIB[4], _3I4551_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_1102_3 (_3I4551_$1I4488_$1I4621_DIB[3], _3I4551_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_1102_2 (_3I4551_$1I4488_$1I4621_DIB[2], _3I4551_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_1102_1 (_3I4551_$1I4488_$1I4621_DIB[1], _3I4551_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_1102_0 (_3I4551_$1I4488_$1I4621_DIB[0], _3I4551_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _3I4551_$1I4488_$1I4621_DIPA;
 reg [1:16] _3I4551_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_1103_0 (_3I4551_$1I4488_$1I4621_DIPA[0], _3I4551_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _3I4551_$1I4488_$1I4621_DIPB;
 reg [1:16] _3I4551_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_1104_1 (_3I4551_$1I4488_$1I4621_DIPB[1], _3I4551_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_1104_0 (_3I4551_$1I4488_$1I4621_DIPB[0], _3I4551_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _3I4551_$1I4488_$1I4621_ENA;
 reg [1:16] _3I4551_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_1105 (_3I4551_$1I4488_$1I4621_ENA, _3I4551_$1I4488_$1I4621_ENA__vlIN);

 wire  _3I4551_$1I4488_$1I4621_ENB;
 reg [1:16] _3I4551_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_1106 (_3I4551_$1I4488_$1I4621_ENB, _3I4551_$1I4488_$1I4621_ENB__vlIN);

 wire  _3I4551_$1I4488_$1I4621_SSRA;
 reg [1:16] _3I4551_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_1107 (_3I4551_$1I4488_$1I4621_SSRA, _3I4551_$1I4488_$1I4621_SSRA__vlIN);

 wire  _3I4551_$1I4488_$1I4621_SSRB;
 reg [1:16] _3I4551_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_1108 (_3I4551_$1I4488_$1I4621_SSRB, _3I4551_$1I4488_$1I4621_SSRB__vlIN);

 wire  _3I4551_$1I4488_$1I4621_WEA;
 reg [1:16] _3I4551_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_1109 (_3I4551_$1I4488_$1I4621_WEA, _3I4551_$1I4488_$1I4621_WEA__vlIN);

 wire  _3I4551_$1I4488_$1I4621_WEB;
 reg [1:16] _3I4551_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_1110 (_3I4551_$1I4488_$1I4621_WEB, _3I4551_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _3I4551_$1I4488_$1I4621 ( _3I4551_$1I4488_$1I4621_DOA , _3I4551_$1I4488_$1I4621_DOB , _3I4551_$1I4488_$1I4621_DOPA , _3I4551_$1I4488_$1I4621_DOPB , _3I4551_$1I4488_$1I4621_ADDRA , _3I4551_$1I4488_$1I4621_ADDRB , _3I4551_$1I4488_$1I4621_CLKA , _3I4551_$1I4488_$1I4621_CLKB , _3I4551_$1I4488_$1I4621_DIA , _3I4551_$1I4488_$1I4621_DIB , _3I4551_$1I4488_$1I4621_DIPA , _3I4551_$1I4488_$1I4621_DIPB , _3I4551_$1I4488_$1I4621_ENA , _3I4551_$1I4488_$1I4621_ENB , _3I4551_$1I4488_$1I4621_SSRA , _3I4551_$1I4488_$1I4621_SSRB , _3I4551_$1I4488_$1I4621_WEA , _3I4551_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4551_$1I4488_$1I4620_DOA;

 wire [15:0] _3I4551_$1I4488_$1I4620_DOB;

 wire [0:0] _3I4551_$1I4488_$1I4620_DOPA;

 wire [1:0] _3I4551_$1I4488_$1I4620_DOPB;

 wire [10:0] _3I4551_$1I4488_$1I4620_ADDRA;
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_1111_10 (_3I4551_$1I4488_$1I4620_ADDRA[10], _3I4551_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_1111_9 (_3I4551_$1I4488_$1I4620_ADDRA[9], _3I4551_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_1111_8 (_3I4551_$1I4488_$1I4620_ADDRA[8], _3I4551_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_1111_7 (_3I4551_$1I4488_$1I4620_ADDRA[7], _3I4551_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_1111_6 (_3I4551_$1I4488_$1I4620_ADDRA[6], _3I4551_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_1111_5 (_3I4551_$1I4488_$1I4620_ADDRA[5], _3I4551_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_1111_4 (_3I4551_$1I4488_$1I4620_ADDRA[4], _3I4551_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_1111_3 (_3I4551_$1I4488_$1I4620_ADDRA[3], _3I4551_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_1111_2 (_3I4551_$1I4488_$1I4620_ADDRA[2], _3I4551_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_1111_1 (_3I4551_$1I4488_$1I4620_ADDRA[1], _3I4551_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_1111_0 (_3I4551_$1I4488_$1I4620_ADDRA[0], _3I4551_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _3I4551_$1I4488_$1I4620_ADDRB;
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1112_9 (_3I4551_$1I4488_$1I4620_ADDRB[9], _3I4551_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1112_8 (_3I4551_$1I4488_$1I4620_ADDRB[8], _3I4551_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1112_7 (_3I4551_$1I4488_$1I4620_ADDRB[7], _3I4551_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1112_6 (_3I4551_$1I4488_$1I4620_ADDRB[6], _3I4551_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1112_5 (_3I4551_$1I4488_$1I4620_ADDRB[5], _3I4551_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1112_4 (_3I4551_$1I4488_$1I4620_ADDRB[4], _3I4551_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1112_3 (_3I4551_$1I4488_$1I4620_ADDRB[3], _3I4551_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1112_2 (_3I4551_$1I4488_$1I4620_ADDRB[2], _3I4551_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1112_1 (_3I4551_$1I4488_$1I4620_ADDRB[1], _3I4551_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1112_0 (_3I4551_$1I4488_$1I4620_ADDRB[0], _3I4551_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _3I4551_$1I4488_$1I4620_CLKA;
 reg [1:16] _3I4551_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1113 (_3I4551_$1I4488_$1I4620_CLKA, _3I4551_$1I4488_$1I4620_CLKA__vlIN);

 wire  _3I4551_$1I4488_$1I4620_CLKB;
 reg [1:16] _3I4551_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1114 (_3I4551_$1I4488_$1I4620_CLKB, _3I4551_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _3I4551_$1I4488_$1I4620_DIA;
 reg [1:16] _3I4551_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1115_7 (_3I4551_$1I4488_$1I4620_DIA[7], _3I4551_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1115_6 (_3I4551_$1I4488_$1I4620_DIA[6], _3I4551_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1115_5 (_3I4551_$1I4488_$1I4620_DIA[5], _3I4551_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1115_4 (_3I4551_$1I4488_$1I4620_DIA[4], _3I4551_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1115_3 (_3I4551_$1I4488_$1I4620_DIA[3], _3I4551_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1115_2 (_3I4551_$1I4488_$1I4620_DIA[2], _3I4551_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1115_1 (_3I4551_$1I4488_$1I4620_DIA[1], _3I4551_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1115_0 (_3I4551_$1I4488_$1I4620_DIA[0], _3I4551_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _3I4551_$1I4488_$1I4620_DIB;
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1116_15 (_3I4551_$1I4488_$1I4620_DIB[15], _3I4551_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1116_14 (_3I4551_$1I4488_$1I4620_DIB[14], _3I4551_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1116_13 (_3I4551_$1I4488_$1I4620_DIB[13], _3I4551_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1116_12 (_3I4551_$1I4488_$1I4620_DIB[12], _3I4551_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1116_11 (_3I4551_$1I4488_$1I4620_DIB[11], _3I4551_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1116_10 (_3I4551_$1I4488_$1I4620_DIB[10], _3I4551_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1116_9 (_3I4551_$1I4488_$1I4620_DIB[9], _3I4551_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1116_8 (_3I4551_$1I4488_$1I4620_DIB[8], _3I4551_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1116_7 (_3I4551_$1I4488_$1I4620_DIB[7], _3I4551_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1116_6 (_3I4551_$1I4488_$1I4620_DIB[6], _3I4551_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1116_5 (_3I4551_$1I4488_$1I4620_DIB[5], _3I4551_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1116_4 (_3I4551_$1I4488_$1I4620_DIB[4], _3I4551_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1116_3 (_3I4551_$1I4488_$1I4620_DIB[3], _3I4551_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1116_2 (_3I4551_$1I4488_$1I4620_DIB[2], _3I4551_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1116_1 (_3I4551_$1I4488_$1I4620_DIB[1], _3I4551_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1116_0 (_3I4551_$1I4488_$1I4620_DIB[0], _3I4551_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _3I4551_$1I4488_$1I4620_DIPA;
 reg [1:16] _3I4551_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1117_0 (_3I4551_$1I4488_$1I4620_DIPA[0], _3I4551_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _3I4551_$1I4488_$1I4620_DIPB;
 reg [1:16] _3I4551_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1118_1 (_3I4551_$1I4488_$1I4620_DIPB[1], _3I4551_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _3I4551_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1118_0 (_3I4551_$1I4488_$1I4620_DIPB[0], _3I4551_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _3I4551_$1I4488_$1I4620_ENA;
 reg [1:16] _3I4551_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1119 (_3I4551_$1I4488_$1I4620_ENA, _3I4551_$1I4488_$1I4620_ENA__vlIN);

 wire  _3I4551_$1I4488_$1I4620_ENB;
 reg [1:16] _3I4551_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1120 (_3I4551_$1I4488_$1I4620_ENB, _3I4551_$1I4488_$1I4620_ENB__vlIN);

 wire  _3I4551_$1I4488_$1I4620_SSRA;
 reg [1:16] _3I4551_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1121 (_3I4551_$1I4488_$1I4620_SSRA, _3I4551_$1I4488_$1I4620_SSRA__vlIN);

 wire  _3I4551_$1I4488_$1I4620_SSRB;
 reg [1:16] _3I4551_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1122 (_3I4551_$1I4488_$1I4620_SSRB, _3I4551_$1I4488_$1I4620_SSRB__vlIN);

 wire  _3I4551_$1I4488_$1I4620_WEA;
 reg [1:16] _3I4551_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1123 (_3I4551_$1I4488_$1I4620_WEA, _3I4551_$1I4488_$1I4620_WEA__vlIN);

 wire  _3I4551_$1I4488_$1I4620_WEB;
 reg [1:16] _3I4551_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1124 (_3I4551_$1I4488_$1I4620_WEB, _3I4551_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _3I4551_$1I4488_$1I4620 ( _3I4551_$1I4488_$1I4620_DOA , _3I4551_$1I4488_$1I4620_DOB , _3I4551_$1I4488_$1I4620_DOPA , _3I4551_$1I4488_$1I4620_DOPB , _3I4551_$1I4488_$1I4620_ADDRA , _3I4551_$1I4488_$1I4620_ADDRB , _3I4551_$1I4488_$1I4620_CLKA , _3I4551_$1I4488_$1I4620_CLKB , _3I4551_$1I4488_$1I4620_DIA , _3I4551_$1I4488_$1I4620_DIB , _3I4551_$1I4488_$1I4620_DIPA , _3I4551_$1I4488_$1I4620_DIPB , _3I4551_$1I4488_$1I4620_ENA , _3I4551_$1I4488_$1I4620_ENB , _3I4551_$1I4488_$1I4620_SSRA , _3I4551_$1I4488_$1I4620_SSRB , _3I4551_$1I4488_$1I4620_WEA , _3I4551_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4526_$1I4488_$1I4621_DOA;

 wire [15:0] _3I4526_$1I4488_$1I4621_DOB;

 wire [0:0] _3I4526_$1I4488_$1I4621_DOPA;

 wire [1:0] _3I4526_$1I4488_$1I4621_DOPB;

 wire [10:0] _3I4526_$1I4488_$1I4621_ADDRA;
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1125_10 (_3I4526_$1I4488_$1I4621_ADDRA[10], _3I4526_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1125_9 (_3I4526_$1I4488_$1I4621_ADDRA[9], _3I4526_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1125_8 (_3I4526_$1I4488_$1I4621_ADDRA[8], _3I4526_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1125_7 (_3I4526_$1I4488_$1I4621_ADDRA[7], _3I4526_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1125_6 (_3I4526_$1I4488_$1I4621_ADDRA[6], _3I4526_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1125_5 (_3I4526_$1I4488_$1I4621_ADDRA[5], _3I4526_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1125_4 (_3I4526_$1I4488_$1I4621_ADDRA[4], _3I4526_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1125_3 (_3I4526_$1I4488_$1I4621_ADDRA[3], _3I4526_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1125_2 (_3I4526_$1I4488_$1I4621_ADDRA[2], _3I4526_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1125_1 (_3I4526_$1I4488_$1I4621_ADDRA[1], _3I4526_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1125_0 (_3I4526_$1I4488_$1I4621_ADDRA[0], _3I4526_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _3I4526_$1I4488_$1I4621_ADDRB;
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_1126_9 (_3I4526_$1I4488_$1I4621_ADDRB[9], _3I4526_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_1126_8 (_3I4526_$1I4488_$1I4621_ADDRB[8], _3I4526_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_1126_7 (_3I4526_$1I4488_$1I4621_ADDRB[7], _3I4526_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_1126_6 (_3I4526_$1I4488_$1I4621_ADDRB[6], _3I4526_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_1126_5 (_3I4526_$1I4488_$1I4621_ADDRB[5], _3I4526_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_1126_4 (_3I4526_$1I4488_$1I4621_ADDRB[4], _3I4526_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_1126_3 (_3I4526_$1I4488_$1I4621_ADDRB[3], _3I4526_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_1126_2 (_3I4526_$1I4488_$1I4621_ADDRB[2], _3I4526_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_1126_1 (_3I4526_$1I4488_$1I4621_ADDRB[1], _3I4526_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_1126_0 (_3I4526_$1I4488_$1I4621_ADDRB[0], _3I4526_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _3I4526_$1I4488_$1I4621_CLKA;
 reg [1:16] _3I4526_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_1127 (_3I4526_$1I4488_$1I4621_CLKA, _3I4526_$1I4488_$1I4621_CLKA__vlIN);

 wire  _3I4526_$1I4488_$1I4621_CLKB;
 reg [1:16] _3I4526_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_1128 (_3I4526_$1I4488_$1I4621_CLKB, _3I4526_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _3I4526_$1I4488_$1I4621_DIA;
 reg [1:16] _3I4526_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_1129_7 (_3I4526_$1I4488_$1I4621_DIA[7], _3I4526_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_1129_6 (_3I4526_$1I4488_$1I4621_DIA[6], _3I4526_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_1129_5 (_3I4526_$1I4488_$1I4621_DIA[5], _3I4526_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_1129_4 (_3I4526_$1I4488_$1I4621_DIA[4], _3I4526_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_1129_3 (_3I4526_$1I4488_$1I4621_DIA[3], _3I4526_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_1129_2 (_3I4526_$1I4488_$1I4621_DIA[2], _3I4526_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_1129_1 (_3I4526_$1I4488_$1I4621_DIA[1], _3I4526_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_1129_0 (_3I4526_$1I4488_$1I4621_DIA[0], _3I4526_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _3I4526_$1I4488_$1I4621_DIB;
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_1130_15 (_3I4526_$1I4488_$1I4621_DIB[15], _3I4526_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_1130_14 (_3I4526_$1I4488_$1I4621_DIB[14], _3I4526_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_1130_13 (_3I4526_$1I4488_$1I4621_DIB[13], _3I4526_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_1130_12 (_3I4526_$1I4488_$1I4621_DIB[12], _3I4526_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_1130_11 (_3I4526_$1I4488_$1I4621_DIB[11], _3I4526_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_1130_10 (_3I4526_$1I4488_$1I4621_DIB[10], _3I4526_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_1130_9 (_3I4526_$1I4488_$1I4621_DIB[9], _3I4526_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_1130_8 (_3I4526_$1I4488_$1I4621_DIB[8], _3I4526_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_1130_7 (_3I4526_$1I4488_$1I4621_DIB[7], _3I4526_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_1130_6 (_3I4526_$1I4488_$1I4621_DIB[6], _3I4526_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_1130_5 (_3I4526_$1I4488_$1I4621_DIB[5], _3I4526_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_1130_4 (_3I4526_$1I4488_$1I4621_DIB[4], _3I4526_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_1130_3 (_3I4526_$1I4488_$1I4621_DIB[3], _3I4526_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_1130_2 (_3I4526_$1I4488_$1I4621_DIB[2], _3I4526_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_1130_1 (_3I4526_$1I4488_$1I4621_DIB[1], _3I4526_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_1130_0 (_3I4526_$1I4488_$1I4621_DIB[0], _3I4526_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _3I4526_$1I4488_$1I4621_DIPA;
 reg [1:16] _3I4526_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_1131_0 (_3I4526_$1I4488_$1I4621_DIPA[0], _3I4526_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _3I4526_$1I4488_$1I4621_DIPB;
 reg [1:16] _3I4526_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_1132_1 (_3I4526_$1I4488_$1I4621_DIPB[1], _3I4526_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_1132_0 (_3I4526_$1I4488_$1I4621_DIPB[0], _3I4526_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _3I4526_$1I4488_$1I4621_ENA;
 reg [1:16] _3I4526_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_1133 (_3I4526_$1I4488_$1I4621_ENA, _3I4526_$1I4488_$1I4621_ENA__vlIN);

 wire  _3I4526_$1I4488_$1I4621_ENB;
 reg [1:16] _3I4526_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_1134 (_3I4526_$1I4488_$1I4621_ENB, _3I4526_$1I4488_$1I4621_ENB__vlIN);

 wire  _3I4526_$1I4488_$1I4621_SSRA;
 reg [1:16] _3I4526_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_1135 (_3I4526_$1I4488_$1I4621_SSRA, _3I4526_$1I4488_$1I4621_SSRA__vlIN);

 wire  _3I4526_$1I4488_$1I4621_SSRB;
 reg [1:16] _3I4526_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_1136 (_3I4526_$1I4488_$1I4621_SSRB, _3I4526_$1I4488_$1I4621_SSRB__vlIN);

 wire  _3I4526_$1I4488_$1I4621_WEA;
 reg [1:16] _3I4526_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_1137 (_3I4526_$1I4488_$1I4621_WEA, _3I4526_$1I4488_$1I4621_WEA__vlIN);

 wire  _3I4526_$1I4488_$1I4621_WEB;
 reg [1:16] _3I4526_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_1138 (_3I4526_$1I4488_$1I4621_WEB, _3I4526_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _3I4526_$1I4488_$1I4621 ( _3I4526_$1I4488_$1I4621_DOA , _3I4526_$1I4488_$1I4621_DOB , _3I4526_$1I4488_$1I4621_DOPA , _3I4526_$1I4488_$1I4621_DOPB , _3I4526_$1I4488_$1I4621_ADDRA , _3I4526_$1I4488_$1I4621_ADDRB , _3I4526_$1I4488_$1I4621_CLKA , _3I4526_$1I4488_$1I4621_CLKB , _3I4526_$1I4488_$1I4621_DIA , _3I4526_$1I4488_$1I4621_DIB , _3I4526_$1I4488_$1I4621_DIPA , _3I4526_$1I4488_$1I4621_DIPB , _3I4526_$1I4488_$1I4621_ENA , _3I4526_$1I4488_$1I4621_ENB , _3I4526_$1I4488_$1I4621_SSRA , _3I4526_$1I4488_$1I4621_SSRB , _3I4526_$1I4488_$1I4621_WEA , _3I4526_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4526_$1I4488_$1I4620_DOA;

 wire [15:0] _3I4526_$1I4488_$1I4620_DOB;

 wire [0:0] _3I4526_$1I4488_$1I4620_DOPA;

 wire [1:0] _3I4526_$1I4488_$1I4620_DOPB;

 wire [10:0] _3I4526_$1I4488_$1I4620_ADDRA;
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_1139_10 (_3I4526_$1I4488_$1I4620_ADDRA[10], _3I4526_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_1139_9 (_3I4526_$1I4488_$1I4620_ADDRA[9], _3I4526_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_1139_8 (_3I4526_$1I4488_$1I4620_ADDRA[8], _3I4526_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_1139_7 (_3I4526_$1I4488_$1I4620_ADDRA[7], _3I4526_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_1139_6 (_3I4526_$1I4488_$1I4620_ADDRA[6], _3I4526_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_1139_5 (_3I4526_$1I4488_$1I4620_ADDRA[5], _3I4526_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_1139_4 (_3I4526_$1I4488_$1I4620_ADDRA[4], _3I4526_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_1139_3 (_3I4526_$1I4488_$1I4620_ADDRA[3], _3I4526_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_1139_2 (_3I4526_$1I4488_$1I4620_ADDRA[2], _3I4526_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_1139_1 (_3I4526_$1I4488_$1I4620_ADDRA[1], _3I4526_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_1139_0 (_3I4526_$1I4488_$1I4620_ADDRA[0], _3I4526_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _3I4526_$1I4488_$1I4620_ADDRB;
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1140_9 (_3I4526_$1I4488_$1I4620_ADDRB[9], _3I4526_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1140_8 (_3I4526_$1I4488_$1I4620_ADDRB[8], _3I4526_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1140_7 (_3I4526_$1I4488_$1I4620_ADDRB[7], _3I4526_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1140_6 (_3I4526_$1I4488_$1I4620_ADDRB[6], _3I4526_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1140_5 (_3I4526_$1I4488_$1I4620_ADDRB[5], _3I4526_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1140_4 (_3I4526_$1I4488_$1I4620_ADDRB[4], _3I4526_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1140_3 (_3I4526_$1I4488_$1I4620_ADDRB[3], _3I4526_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1140_2 (_3I4526_$1I4488_$1I4620_ADDRB[2], _3I4526_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1140_1 (_3I4526_$1I4488_$1I4620_ADDRB[1], _3I4526_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1140_0 (_3I4526_$1I4488_$1I4620_ADDRB[0], _3I4526_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _3I4526_$1I4488_$1I4620_CLKA;
 reg [1:16] _3I4526_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1141 (_3I4526_$1I4488_$1I4620_CLKA, _3I4526_$1I4488_$1I4620_CLKA__vlIN);

 wire  _3I4526_$1I4488_$1I4620_CLKB;
 reg [1:16] _3I4526_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1142 (_3I4526_$1I4488_$1I4620_CLKB, _3I4526_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _3I4526_$1I4488_$1I4620_DIA;
 reg [1:16] _3I4526_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1143_7 (_3I4526_$1I4488_$1I4620_DIA[7], _3I4526_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1143_6 (_3I4526_$1I4488_$1I4620_DIA[6], _3I4526_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1143_5 (_3I4526_$1I4488_$1I4620_DIA[5], _3I4526_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1143_4 (_3I4526_$1I4488_$1I4620_DIA[4], _3I4526_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1143_3 (_3I4526_$1I4488_$1I4620_DIA[3], _3I4526_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1143_2 (_3I4526_$1I4488_$1I4620_DIA[2], _3I4526_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1143_1 (_3I4526_$1I4488_$1I4620_DIA[1], _3I4526_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1143_0 (_3I4526_$1I4488_$1I4620_DIA[0], _3I4526_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _3I4526_$1I4488_$1I4620_DIB;
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1144_15 (_3I4526_$1I4488_$1I4620_DIB[15], _3I4526_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1144_14 (_3I4526_$1I4488_$1I4620_DIB[14], _3I4526_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1144_13 (_3I4526_$1I4488_$1I4620_DIB[13], _3I4526_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1144_12 (_3I4526_$1I4488_$1I4620_DIB[12], _3I4526_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1144_11 (_3I4526_$1I4488_$1I4620_DIB[11], _3I4526_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1144_10 (_3I4526_$1I4488_$1I4620_DIB[10], _3I4526_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1144_9 (_3I4526_$1I4488_$1I4620_DIB[9], _3I4526_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1144_8 (_3I4526_$1I4488_$1I4620_DIB[8], _3I4526_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1144_7 (_3I4526_$1I4488_$1I4620_DIB[7], _3I4526_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1144_6 (_3I4526_$1I4488_$1I4620_DIB[6], _3I4526_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1144_5 (_3I4526_$1I4488_$1I4620_DIB[5], _3I4526_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1144_4 (_3I4526_$1I4488_$1I4620_DIB[4], _3I4526_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1144_3 (_3I4526_$1I4488_$1I4620_DIB[3], _3I4526_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1144_2 (_3I4526_$1I4488_$1I4620_DIB[2], _3I4526_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1144_1 (_3I4526_$1I4488_$1I4620_DIB[1], _3I4526_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1144_0 (_3I4526_$1I4488_$1I4620_DIB[0], _3I4526_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _3I4526_$1I4488_$1I4620_DIPA;
 reg [1:16] _3I4526_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1145_0 (_3I4526_$1I4488_$1I4620_DIPA[0], _3I4526_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _3I4526_$1I4488_$1I4620_DIPB;
 reg [1:16] _3I4526_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1146_1 (_3I4526_$1I4488_$1I4620_DIPB[1], _3I4526_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _3I4526_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1146_0 (_3I4526_$1I4488_$1I4620_DIPB[0], _3I4526_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _3I4526_$1I4488_$1I4620_ENA;
 reg [1:16] _3I4526_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1147 (_3I4526_$1I4488_$1I4620_ENA, _3I4526_$1I4488_$1I4620_ENA__vlIN);

 wire  _3I4526_$1I4488_$1I4620_ENB;
 reg [1:16] _3I4526_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1148 (_3I4526_$1I4488_$1I4620_ENB, _3I4526_$1I4488_$1I4620_ENB__vlIN);

 wire  _3I4526_$1I4488_$1I4620_SSRA;
 reg [1:16] _3I4526_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1149 (_3I4526_$1I4488_$1I4620_SSRA, _3I4526_$1I4488_$1I4620_SSRA__vlIN);

 wire  _3I4526_$1I4488_$1I4620_SSRB;
 reg [1:16] _3I4526_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1150 (_3I4526_$1I4488_$1I4620_SSRB, _3I4526_$1I4488_$1I4620_SSRB__vlIN);

 wire  _3I4526_$1I4488_$1I4620_WEA;
 reg [1:16] _3I4526_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1151 (_3I4526_$1I4488_$1I4620_WEA, _3I4526_$1I4488_$1I4620_WEA__vlIN);

 wire  _3I4526_$1I4488_$1I4620_WEB;
 reg [1:16] _3I4526_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1152 (_3I4526_$1I4488_$1I4620_WEB, _3I4526_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _3I4526_$1I4488_$1I4620 ( _3I4526_$1I4488_$1I4620_DOA , _3I4526_$1I4488_$1I4620_DOB , _3I4526_$1I4488_$1I4620_DOPA , _3I4526_$1I4488_$1I4620_DOPB , _3I4526_$1I4488_$1I4620_ADDRA , _3I4526_$1I4488_$1I4620_ADDRB , _3I4526_$1I4488_$1I4620_CLKA , _3I4526_$1I4488_$1I4620_CLKB , _3I4526_$1I4488_$1I4620_DIA , _3I4526_$1I4488_$1I4620_DIB , _3I4526_$1I4488_$1I4620_DIPA , _3I4526_$1I4488_$1I4620_DIPB , _3I4526_$1I4488_$1I4620_ENA , _3I4526_$1I4488_$1I4620_ENB , _3I4526_$1I4488_$1I4620_SSRA , _3I4526_$1I4488_$1I4620_SSRB , _3I4526_$1I4488_$1I4620_WEA , _3I4526_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4496_$1I4488_$1I4621_DOA;

 wire [15:0] _3I4496_$1I4488_$1I4621_DOB;

 wire [0:0] _3I4496_$1I4488_$1I4621_DOPA;

 wire [1:0] _3I4496_$1I4488_$1I4621_DOPB;

 wire [10:0] _3I4496_$1I4488_$1I4621_ADDRA;
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1153_10 (_3I4496_$1I4488_$1I4621_ADDRA[10], _3I4496_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1153_9 (_3I4496_$1I4488_$1I4621_ADDRA[9], _3I4496_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1153_8 (_3I4496_$1I4488_$1I4621_ADDRA[8], _3I4496_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1153_7 (_3I4496_$1I4488_$1I4621_ADDRA[7], _3I4496_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1153_6 (_3I4496_$1I4488_$1I4621_ADDRA[6], _3I4496_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1153_5 (_3I4496_$1I4488_$1I4621_ADDRA[5], _3I4496_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1153_4 (_3I4496_$1I4488_$1I4621_ADDRA[4], _3I4496_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1153_3 (_3I4496_$1I4488_$1I4621_ADDRA[3], _3I4496_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1153_2 (_3I4496_$1I4488_$1I4621_ADDRA[2], _3I4496_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1153_1 (_3I4496_$1I4488_$1I4621_ADDRA[1], _3I4496_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1153_0 (_3I4496_$1I4488_$1I4621_ADDRA[0], _3I4496_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _3I4496_$1I4488_$1I4621_ADDRB;
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_1154_9 (_3I4496_$1I4488_$1I4621_ADDRB[9], _3I4496_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_1154_8 (_3I4496_$1I4488_$1I4621_ADDRB[8], _3I4496_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_1154_7 (_3I4496_$1I4488_$1I4621_ADDRB[7], _3I4496_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_1154_6 (_3I4496_$1I4488_$1I4621_ADDRB[6], _3I4496_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_1154_5 (_3I4496_$1I4488_$1I4621_ADDRB[5], _3I4496_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_1154_4 (_3I4496_$1I4488_$1I4621_ADDRB[4], _3I4496_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_1154_3 (_3I4496_$1I4488_$1I4621_ADDRB[3], _3I4496_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_1154_2 (_3I4496_$1I4488_$1I4621_ADDRB[2], _3I4496_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_1154_1 (_3I4496_$1I4488_$1I4621_ADDRB[1], _3I4496_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_1154_0 (_3I4496_$1I4488_$1I4621_ADDRB[0], _3I4496_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _3I4496_$1I4488_$1I4621_CLKA;
 reg [1:16] _3I4496_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_1155 (_3I4496_$1I4488_$1I4621_CLKA, _3I4496_$1I4488_$1I4621_CLKA__vlIN);

 wire  _3I4496_$1I4488_$1I4621_CLKB;
 reg [1:16] _3I4496_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_1156 (_3I4496_$1I4488_$1I4621_CLKB, _3I4496_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _3I4496_$1I4488_$1I4621_DIA;
 reg [1:16] _3I4496_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_1157_7 (_3I4496_$1I4488_$1I4621_DIA[7], _3I4496_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_1157_6 (_3I4496_$1I4488_$1I4621_DIA[6], _3I4496_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_1157_5 (_3I4496_$1I4488_$1I4621_DIA[5], _3I4496_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_1157_4 (_3I4496_$1I4488_$1I4621_DIA[4], _3I4496_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_1157_3 (_3I4496_$1I4488_$1I4621_DIA[3], _3I4496_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_1157_2 (_3I4496_$1I4488_$1I4621_DIA[2], _3I4496_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_1157_1 (_3I4496_$1I4488_$1I4621_DIA[1], _3I4496_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_1157_0 (_3I4496_$1I4488_$1I4621_DIA[0], _3I4496_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _3I4496_$1I4488_$1I4621_DIB;
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_1158_15 (_3I4496_$1I4488_$1I4621_DIB[15], _3I4496_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_1158_14 (_3I4496_$1I4488_$1I4621_DIB[14], _3I4496_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_1158_13 (_3I4496_$1I4488_$1I4621_DIB[13], _3I4496_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_1158_12 (_3I4496_$1I4488_$1I4621_DIB[12], _3I4496_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_1158_11 (_3I4496_$1I4488_$1I4621_DIB[11], _3I4496_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_1158_10 (_3I4496_$1I4488_$1I4621_DIB[10], _3I4496_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_1158_9 (_3I4496_$1I4488_$1I4621_DIB[9], _3I4496_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_1158_8 (_3I4496_$1I4488_$1I4621_DIB[8], _3I4496_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_1158_7 (_3I4496_$1I4488_$1I4621_DIB[7], _3I4496_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_1158_6 (_3I4496_$1I4488_$1I4621_DIB[6], _3I4496_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_1158_5 (_3I4496_$1I4488_$1I4621_DIB[5], _3I4496_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_1158_4 (_3I4496_$1I4488_$1I4621_DIB[4], _3I4496_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_1158_3 (_3I4496_$1I4488_$1I4621_DIB[3], _3I4496_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_1158_2 (_3I4496_$1I4488_$1I4621_DIB[2], _3I4496_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_1158_1 (_3I4496_$1I4488_$1I4621_DIB[1], _3I4496_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_1158_0 (_3I4496_$1I4488_$1I4621_DIB[0], _3I4496_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _3I4496_$1I4488_$1I4621_DIPA;
 reg [1:16] _3I4496_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_1159_0 (_3I4496_$1I4488_$1I4621_DIPA[0], _3I4496_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _3I4496_$1I4488_$1I4621_DIPB;
 reg [1:16] _3I4496_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_1160_1 (_3I4496_$1I4488_$1I4621_DIPB[1], _3I4496_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_1160_0 (_3I4496_$1I4488_$1I4621_DIPB[0], _3I4496_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _3I4496_$1I4488_$1I4621_ENA;
 reg [1:16] _3I4496_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_1161 (_3I4496_$1I4488_$1I4621_ENA, _3I4496_$1I4488_$1I4621_ENA__vlIN);

 wire  _3I4496_$1I4488_$1I4621_ENB;
 reg [1:16] _3I4496_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_1162 (_3I4496_$1I4488_$1I4621_ENB, _3I4496_$1I4488_$1I4621_ENB__vlIN);

 wire  _3I4496_$1I4488_$1I4621_SSRA;
 reg [1:16] _3I4496_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_1163 (_3I4496_$1I4488_$1I4621_SSRA, _3I4496_$1I4488_$1I4621_SSRA__vlIN);

 wire  _3I4496_$1I4488_$1I4621_SSRB;
 reg [1:16] _3I4496_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_1164 (_3I4496_$1I4488_$1I4621_SSRB, _3I4496_$1I4488_$1I4621_SSRB__vlIN);

 wire  _3I4496_$1I4488_$1I4621_WEA;
 reg [1:16] _3I4496_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_1165 (_3I4496_$1I4488_$1I4621_WEA, _3I4496_$1I4488_$1I4621_WEA__vlIN);

 wire  _3I4496_$1I4488_$1I4621_WEB;
 reg [1:16] _3I4496_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_1166 (_3I4496_$1I4488_$1I4621_WEB, _3I4496_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _3I4496_$1I4488_$1I4621 ( _3I4496_$1I4488_$1I4621_DOA , _3I4496_$1I4488_$1I4621_DOB , _3I4496_$1I4488_$1I4621_DOPA , _3I4496_$1I4488_$1I4621_DOPB , _3I4496_$1I4488_$1I4621_ADDRA , _3I4496_$1I4488_$1I4621_ADDRB , _3I4496_$1I4488_$1I4621_CLKA , _3I4496_$1I4488_$1I4621_CLKB , _3I4496_$1I4488_$1I4621_DIA , _3I4496_$1I4488_$1I4621_DIB , _3I4496_$1I4488_$1I4621_DIPA , _3I4496_$1I4488_$1I4621_DIPB , _3I4496_$1I4488_$1I4621_ENA , _3I4496_$1I4488_$1I4621_ENB , _3I4496_$1I4488_$1I4621_SSRA , _3I4496_$1I4488_$1I4621_SSRB , _3I4496_$1I4488_$1I4621_WEA , _3I4496_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4496_$1I4488_$1I4620_DOA;

 wire [15:0] _3I4496_$1I4488_$1I4620_DOB;

 wire [0:0] _3I4496_$1I4488_$1I4620_DOPA;

 wire [1:0] _3I4496_$1I4488_$1I4620_DOPB;

 wire [10:0] _3I4496_$1I4488_$1I4620_ADDRA;
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_1167_10 (_3I4496_$1I4488_$1I4620_ADDRA[10], _3I4496_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_1167_9 (_3I4496_$1I4488_$1I4620_ADDRA[9], _3I4496_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_1167_8 (_3I4496_$1I4488_$1I4620_ADDRA[8], _3I4496_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_1167_7 (_3I4496_$1I4488_$1I4620_ADDRA[7], _3I4496_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_1167_6 (_3I4496_$1I4488_$1I4620_ADDRA[6], _3I4496_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_1167_5 (_3I4496_$1I4488_$1I4620_ADDRA[5], _3I4496_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_1167_4 (_3I4496_$1I4488_$1I4620_ADDRA[4], _3I4496_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_1167_3 (_3I4496_$1I4488_$1I4620_ADDRA[3], _3I4496_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_1167_2 (_3I4496_$1I4488_$1I4620_ADDRA[2], _3I4496_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_1167_1 (_3I4496_$1I4488_$1I4620_ADDRA[1], _3I4496_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_1167_0 (_3I4496_$1I4488_$1I4620_ADDRA[0], _3I4496_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _3I4496_$1I4488_$1I4620_ADDRB;
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1168_9 (_3I4496_$1I4488_$1I4620_ADDRB[9], _3I4496_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1168_8 (_3I4496_$1I4488_$1I4620_ADDRB[8], _3I4496_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1168_7 (_3I4496_$1I4488_$1I4620_ADDRB[7], _3I4496_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1168_6 (_3I4496_$1I4488_$1I4620_ADDRB[6], _3I4496_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1168_5 (_3I4496_$1I4488_$1I4620_ADDRB[5], _3I4496_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1168_4 (_3I4496_$1I4488_$1I4620_ADDRB[4], _3I4496_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1168_3 (_3I4496_$1I4488_$1I4620_ADDRB[3], _3I4496_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1168_2 (_3I4496_$1I4488_$1I4620_ADDRB[2], _3I4496_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1168_1 (_3I4496_$1I4488_$1I4620_ADDRB[1], _3I4496_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1168_0 (_3I4496_$1I4488_$1I4620_ADDRB[0], _3I4496_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _3I4496_$1I4488_$1I4620_CLKA;
 reg [1:16] _3I4496_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1169 (_3I4496_$1I4488_$1I4620_CLKA, _3I4496_$1I4488_$1I4620_CLKA__vlIN);

 wire  _3I4496_$1I4488_$1I4620_CLKB;
 reg [1:16] _3I4496_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1170 (_3I4496_$1I4488_$1I4620_CLKB, _3I4496_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _3I4496_$1I4488_$1I4620_DIA;
 reg [1:16] _3I4496_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1171_7 (_3I4496_$1I4488_$1I4620_DIA[7], _3I4496_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1171_6 (_3I4496_$1I4488_$1I4620_DIA[6], _3I4496_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1171_5 (_3I4496_$1I4488_$1I4620_DIA[5], _3I4496_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1171_4 (_3I4496_$1I4488_$1I4620_DIA[4], _3I4496_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1171_3 (_3I4496_$1I4488_$1I4620_DIA[3], _3I4496_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1171_2 (_3I4496_$1I4488_$1I4620_DIA[2], _3I4496_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1171_1 (_3I4496_$1I4488_$1I4620_DIA[1], _3I4496_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1171_0 (_3I4496_$1I4488_$1I4620_DIA[0], _3I4496_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _3I4496_$1I4488_$1I4620_DIB;
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1172_15 (_3I4496_$1I4488_$1I4620_DIB[15], _3I4496_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1172_14 (_3I4496_$1I4488_$1I4620_DIB[14], _3I4496_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1172_13 (_3I4496_$1I4488_$1I4620_DIB[13], _3I4496_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1172_12 (_3I4496_$1I4488_$1I4620_DIB[12], _3I4496_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1172_11 (_3I4496_$1I4488_$1I4620_DIB[11], _3I4496_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1172_10 (_3I4496_$1I4488_$1I4620_DIB[10], _3I4496_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1172_9 (_3I4496_$1I4488_$1I4620_DIB[9], _3I4496_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1172_8 (_3I4496_$1I4488_$1I4620_DIB[8], _3I4496_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1172_7 (_3I4496_$1I4488_$1I4620_DIB[7], _3I4496_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1172_6 (_3I4496_$1I4488_$1I4620_DIB[6], _3I4496_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1172_5 (_3I4496_$1I4488_$1I4620_DIB[5], _3I4496_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1172_4 (_3I4496_$1I4488_$1I4620_DIB[4], _3I4496_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1172_3 (_3I4496_$1I4488_$1I4620_DIB[3], _3I4496_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1172_2 (_3I4496_$1I4488_$1I4620_DIB[2], _3I4496_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1172_1 (_3I4496_$1I4488_$1I4620_DIB[1], _3I4496_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1172_0 (_3I4496_$1I4488_$1I4620_DIB[0], _3I4496_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _3I4496_$1I4488_$1I4620_DIPA;
 reg [1:16] _3I4496_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1173_0 (_3I4496_$1I4488_$1I4620_DIPA[0], _3I4496_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _3I4496_$1I4488_$1I4620_DIPB;
 reg [1:16] _3I4496_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1174_1 (_3I4496_$1I4488_$1I4620_DIPB[1], _3I4496_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _3I4496_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1174_0 (_3I4496_$1I4488_$1I4620_DIPB[0], _3I4496_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _3I4496_$1I4488_$1I4620_ENA;
 reg [1:16] _3I4496_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1175 (_3I4496_$1I4488_$1I4620_ENA, _3I4496_$1I4488_$1I4620_ENA__vlIN);

 wire  _3I4496_$1I4488_$1I4620_ENB;
 reg [1:16] _3I4496_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1176 (_3I4496_$1I4488_$1I4620_ENB, _3I4496_$1I4488_$1I4620_ENB__vlIN);

 wire  _3I4496_$1I4488_$1I4620_SSRA;
 reg [1:16] _3I4496_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1177 (_3I4496_$1I4488_$1I4620_SSRA, _3I4496_$1I4488_$1I4620_SSRA__vlIN);

 wire  _3I4496_$1I4488_$1I4620_SSRB;
 reg [1:16] _3I4496_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1178 (_3I4496_$1I4488_$1I4620_SSRB, _3I4496_$1I4488_$1I4620_SSRB__vlIN);

 wire  _3I4496_$1I4488_$1I4620_WEA;
 reg [1:16] _3I4496_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1179 (_3I4496_$1I4488_$1I4620_WEA, _3I4496_$1I4488_$1I4620_WEA__vlIN);

 wire  _3I4496_$1I4488_$1I4620_WEB;
 reg [1:16] _3I4496_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1180 (_3I4496_$1I4488_$1I4620_WEB, _3I4496_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _3I4496_$1I4488_$1I4620 ( _3I4496_$1I4488_$1I4620_DOA , _3I4496_$1I4488_$1I4620_DOB , _3I4496_$1I4488_$1I4620_DOPA , _3I4496_$1I4488_$1I4620_DOPB , _3I4496_$1I4488_$1I4620_ADDRA , _3I4496_$1I4488_$1I4620_ADDRB , _3I4496_$1I4488_$1I4620_CLKA , _3I4496_$1I4488_$1I4620_CLKB , _3I4496_$1I4488_$1I4620_DIA , _3I4496_$1I4488_$1I4620_DIB , _3I4496_$1I4488_$1I4620_DIPA , _3I4496_$1I4488_$1I4620_DIPB , _3I4496_$1I4488_$1I4620_ENA , _3I4496_$1I4488_$1I4620_ENB , _3I4496_$1I4488_$1I4620_SSRA , _3I4496_$1I4488_$1I4620_SSRB , _3I4496_$1I4488_$1I4620_WEA , _3I4496_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4489_$1I4488_$1I4621_DOA;

 wire [15:0] _3I4489_$1I4488_$1I4621_DOB;

 wire [0:0] _3I4489_$1I4488_$1I4621_DOPA;

 wire [1:0] _3I4489_$1I4488_$1I4621_DOPB;

 wire [10:0] _3I4489_$1I4488_$1I4621_ADDRA;
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1181_10 (_3I4489_$1I4488_$1I4621_ADDRA[10], _3I4489_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1181_9 (_3I4489_$1I4488_$1I4621_ADDRA[9], _3I4489_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1181_8 (_3I4489_$1I4488_$1I4621_ADDRA[8], _3I4489_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1181_7 (_3I4489_$1I4488_$1I4621_ADDRA[7], _3I4489_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1181_6 (_3I4489_$1I4488_$1I4621_ADDRA[6], _3I4489_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1181_5 (_3I4489_$1I4488_$1I4621_ADDRA[5], _3I4489_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1181_4 (_3I4489_$1I4488_$1I4621_ADDRA[4], _3I4489_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1181_3 (_3I4489_$1I4488_$1I4621_ADDRA[3], _3I4489_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1181_2 (_3I4489_$1I4488_$1I4621_ADDRA[2], _3I4489_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1181_1 (_3I4489_$1I4488_$1I4621_ADDRA[1], _3I4489_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1181_0 (_3I4489_$1I4488_$1I4621_ADDRA[0], _3I4489_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _3I4489_$1I4488_$1I4621_ADDRB;
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_1182_9 (_3I4489_$1I4488_$1I4621_ADDRB[9], _3I4489_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_1182_8 (_3I4489_$1I4488_$1I4621_ADDRB[8], _3I4489_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_1182_7 (_3I4489_$1I4488_$1I4621_ADDRB[7], _3I4489_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_1182_6 (_3I4489_$1I4488_$1I4621_ADDRB[6], _3I4489_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_1182_5 (_3I4489_$1I4488_$1I4621_ADDRB[5], _3I4489_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_1182_4 (_3I4489_$1I4488_$1I4621_ADDRB[4], _3I4489_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_1182_3 (_3I4489_$1I4488_$1I4621_ADDRB[3], _3I4489_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_1182_2 (_3I4489_$1I4488_$1I4621_ADDRB[2], _3I4489_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_1182_1 (_3I4489_$1I4488_$1I4621_ADDRB[1], _3I4489_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_1182_0 (_3I4489_$1I4488_$1I4621_ADDRB[0], _3I4489_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _3I4489_$1I4488_$1I4621_CLKA;
 reg [1:16] _3I4489_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_1183 (_3I4489_$1I4488_$1I4621_CLKA, _3I4489_$1I4488_$1I4621_CLKA__vlIN);

 wire  _3I4489_$1I4488_$1I4621_CLKB;
 reg [1:16] _3I4489_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_1184 (_3I4489_$1I4488_$1I4621_CLKB, _3I4489_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _3I4489_$1I4488_$1I4621_DIA;
 reg [1:16] _3I4489_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_1185_7 (_3I4489_$1I4488_$1I4621_DIA[7], _3I4489_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_1185_6 (_3I4489_$1I4488_$1I4621_DIA[6], _3I4489_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_1185_5 (_3I4489_$1I4488_$1I4621_DIA[5], _3I4489_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_1185_4 (_3I4489_$1I4488_$1I4621_DIA[4], _3I4489_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_1185_3 (_3I4489_$1I4488_$1I4621_DIA[3], _3I4489_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_1185_2 (_3I4489_$1I4488_$1I4621_DIA[2], _3I4489_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_1185_1 (_3I4489_$1I4488_$1I4621_DIA[1], _3I4489_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_1185_0 (_3I4489_$1I4488_$1I4621_DIA[0], _3I4489_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _3I4489_$1I4488_$1I4621_DIB;
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_1186_15 (_3I4489_$1I4488_$1I4621_DIB[15], _3I4489_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_1186_14 (_3I4489_$1I4488_$1I4621_DIB[14], _3I4489_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_1186_13 (_3I4489_$1I4488_$1I4621_DIB[13], _3I4489_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_1186_12 (_3I4489_$1I4488_$1I4621_DIB[12], _3I4489_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_1186_11 (_3I4489_$1I4488_$1I4621_DIB[11], _3I4489_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_1186_10 (_3I4489_$1I4488_$1I4621_DIB[10], _3I4489_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_1186_9 (_3I4489_$1I4488_$1I4621_DIB[9], _3I4489_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_1186_8 (_3I4489_$1I4488_$1I4621_DIB[8], _3I4489_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_1186_7 (_3I4489_$1I4488_$1I4621_DIB[7], _3I4489_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_1186_6 (_3I4489_$1I4488_$1I4621_DIB[6], _3I4489_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_1186_5 (_3I4489_$1I4488_$1I4621_DIB[5], _3I4489_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_1186_4 (_3I4489_$1I4488_$1I4621_DIB[4], _3I4489_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_1186_3 (_3I4489_$1I4488_$1I4621_DIB[3], _3I4489_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_1186_2 (_3I4489_$1I4488_$1I4621_DIB[2], _3I4489_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_1186_1 (_3I4489_$1I4488_$1I4621_DIB[1], _3I4489_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_1186_0 (_3I4489_$1I4488_$1I4621_DIB[0], _3I4489_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _3I4489_$1I4488_$1I4621_DIPA;
 reg [1:16] _3I4489_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_1187_0 (_3I4489_$1I4488_$1I4621_DIPA[0], _3I4489_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _3I4489_$1I4488_$1I4621_DIPB;
 reg [1:16] _3I4489_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_1188_1 (_3I4489_$1I4488_$1I4621_DIPB[1], _3I4489_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_1188_0 (_3I4489_$1I4488_$1I4621_DIPB[0], _3I4489_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _3I4489_$1I4488_$1I4621_ENA;
 reg [1:16] _3I4489_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_1189 (_3I4489_$1I4488_$1I4621_ENA, _3I4489_$1I4488_$1I4621_ENA__vlIN);

 wire  _3I4489_$1I4488_$1I4621_ENB;
 reg [1:16] _3I4489_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_1190 (_3I4489_$1I4488_$1I4621_ENB, _3I4489_$1I4488_$1I4621_ENB__vlIN);

 wire  _3I4489_$1I4488_$1I4621_SSRA;
 reg [1:16] _3I4489_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_1191 (_3I4489_$1I4488_$1I4621_SSRA, _3I4489_$1I4488_$1I4621_SSRA__vlIN);

 wire  _3I4489_$1I4488_$1I4621_SSRB;
 reg [1:16] _3I4489_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_1192 (_3I4489_$1I4488_$1I4621_SSRB, _3I4489_$1I4488_$1I4621_SSRB__vlIN);

 wire  _3I4489_$1I4488_$1I4621_WEA;
 reg [1:16] _3I4489_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_1193 (_3I4489_$1I4488_$1I4621_WEA, _3I4489_$1I4488_$1I4621_WEA__vlIN);

 wire  _3I4489_$1I4488_$1I4621_WEB;
 reg [1:16] _3I4489_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_1194 (_3I4489_$1I4488_$1I4621_WEB, _3I4489_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _3I4489_$1I4488_$1I4621 ( _3I4489_$1I4488_$1I4621_DOA , _3I4489_$1I4488_$1I4621_DOB , _3I4489_$1I4488_$1I4621_DOPA , _3I4489_$1I4488_$1I4621_DOPB , _3I4489_$1I4488_$1I4621_ADDRA , _3I4489_$1I4488_$1I4621_ADDRB , _3I4489_$1I4488_$1I4621_CLKA , _3I4489_$1I4488_$1I4621_CLKB , _3I4489_$1I4488_$1I4621_DIA , _3I4489_$1I4488_$1I4621_DIB , _3I4489_$1I4488_$1I4621_DIPA , _3I4489_$1I4488_$1I4621_DIPB , _3I4489_$1I4488_$1I4621_ENA , _3I4489_$1I4488_$1I4621_ENB , _3I4489_$1I4488_$1I4621_SSRA , _3I4489_$1I4488_$1I4621_SSRB , _3I4489_$1I4488_$1I4621_WEA , _3I4489_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4489_$1I4488_$1I4620_DOA;

 wire [15:0] _3I4489_$1I4488_$1I4620_DOB;

 wire [0:0] _3I4489_$1I4488_$1I4620_DOPA;

 wire [1:0] _3I4489_$1I4488_$1I4620_DOPB;

 wire [10:0] _3I4489_$1I4488_$1I4620_ADDRA;
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_1195_10 (_3I4489_$1I4488_$1I4620_ADDRA[10], _3I4489_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_1195_9 (_3I4489_$1I4488_$1I4620_ADDRA[9], _3I4489_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_1195_8 (_3I4489_$1I4488_$1I4620_ADDRA[8], _3I4489_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_1195_7 (_3I4489_$1I4488_$1I4620_ADDRA[7], _3I4489_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_1195_6 (_3I4489_$1I4488_$1I4620_ADDRA[6], _3I4489_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_1195_5 (_3I4489_$1I4488_$1I4620_ADDRA[5], _3I4489_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_1195_4 (_3I4489_$1I4488_$1I4620_ADDRA[4], _3I4489_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_1195_3 (_3I4489_$1I4488_$1I4620_ADDRA[3], _3I4489_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_1195_2 (_3I4489_$1I4488_$1I4620_ADDRA[2], _3I4489_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_1195_1 (_3I4489_$1I4488_$1I4620_ADDRA[1], _3I4489_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_1195_0 (_3I4489_$1I4488_$1I4620_ADDRA[0], _3I4489_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _3I4489_$1I4488_$1I4620_ADDRB;
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1196_9 (_3I4489_$1I4488_$1I4620_ADDRB[9], _3I4489_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1196_8 (_3I4489_$1I4488_$1I4620_ADDRB[8], _3I4489_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1196_7 (_3I4489_$1I4488_$1I4620_ADDRB[7], _3I4489_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1196_6 (_3I4489_$1I4488_$1I4620_ADDRB[6], _3I4489_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1196_5 (_3I4489_$1I4488_$1I4620_ADDRB[5], _3I4489_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1196_4 (_3I4489_$1I4488_$1I4620_ADDRB[4], _3I4489_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1196_3 (_3I4489_$1I4488_$1I4620_ADDRB[3], _3I4489_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1196_2 (_3I4489_$1I4488_$1I4620_ADDRB[2], _3I4489_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1196_1 (_3I4489_$1I4488_$1I4620_ADDRB[1], _3I4489_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1196_0 (_3I4489_$1I4488_$1I4620_ADDRB[0], _3I4489_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _3I4489_$1I4488_$1I4620_CLKA;
 reg [1:16] _3I4489_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1197 (_3I4489_$1I4488_$1I4620_CLKA, _3I4489_$1I4488_$1I4620_CLKA__vlIN);

 wire  _3I4489_$1I4488_$1I4620_CLKB;
 reg [1:16] _3I4489_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1198 (_3I4489_$1I4488_$1I4620_CLKB, _3I4489_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _3I4489_$1I4488_$1I4620_DIA;
 reg [1:16] _3I4489_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1199_7 (_3I4489_$1I4488_$1I4620_DIA[7], _3I4489_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1199_6 (_3I4489_$1I4488_$1I4620_DIA[6], _3I4489_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1199_5 (_3I4489_$1I4488_$1I4620_DIA[5], _3I4489_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1199_4 (_3I4489_$1I4488_$1I4620_DIA[4], _3I4489_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1199_3 (_3I4489_$1I4488_$1I4620_DIA[3], _3I4489_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1199_2 (_3I4489_$1I4488_$1I4620_DIA[2], _3I4489_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1199_1 (_3I4489_$1I4488_$1I4620_DIA[1], _3I4489_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1199_0 (_3I4489_$1I4488_$1I4620_DIA[0], _3I4489_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _3I4489_$1I4488_$1I4620_DIB;
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1200_15 (_3I4489_$1I4488_$1I4620_DIB[15], _3I4489_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1200_14 (_3I4489_$1I4488_$1I4620_DIB[14], _3I4489_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1200_13 (_3I4489_$1I4488_$1I4620_DIB[13], _3I4489_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1200_12 (_3I4489_$1I4488_$1I4620_DIB[12], _3I4489_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1200_11 (_3I4489_$1I4488_$1I4620_DIB[11], _3I4489_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1200_10 (_3I4489_$1I4488_$1I4620_DIB[10], _3I4489_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1200_9 (_3I4489_$1I4488_$1I4620_DIB[9], _3I4489_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1200_8 (_3I4489_$1I4488_$1I4620_DIB[8], _3I4489_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1200_7 (_3I4489_$1I4488_$1I4620_DIB[7], _3I4489_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1200_6 (_3I4489_$1I4488_$1I4620_DIB[6], _3I4489_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1200_5 (_3I4489_$1I4488_$1I4620_DIB[5], _3I4489_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1200_4 (_3I4489_$1I4488_$1I4620_DIB[4], _3I4489_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1200_3 (_3I4489_$1I4488_$1I4620_DIB[3], _3I4489_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1200_2 (_3I4489_$1I4488_$1I4620_DIB[2], _3I4489_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1200_1 (_3I4489_$1I4488_$1I4620_DIB[1], _3I4489_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1200_0 (_3I4489_$1I4488_$1I4620_DIB[0], _3I4489_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _3I4489_$1I4488_$1I4620_DIPA;
 reg [1:16] _3I4489_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1201_0 (_3I4489_$1I4488_$1I4620_DIPA[0], _3I4489_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _3I4489_$1I4488_$1I4620_DIPB;
 reg [1:16] _3I4489_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1202_1 (_3I4489_$1I4488_$1I4620_DIPB[1], _3I4489_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _3I4489_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1202_0 (_3I4489_$1I4488_$1I4620_DIPB[0], _3I4489_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _3I4489_$1I4488_$1I4620_ENA;
 reg [1:16] _3I4489_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1203 (_3I4489_$1I4488_$1I4620_ENA, _3I4489_$1I4488_$1I4620_ENA__vlIN);

 wire  _3I4489_$1I4488_$1I4620_ENB;
 reg [1:16] _3I4489_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1204 (_3I4489_$1I4488_$1I4620_ENB, _3I4489_$1I4488_$1I4620_ENB__vlIN);

 wire  _3I4489_$1I4488_$1I4620_SSRA;
 reg [1:16] _3I4489_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1205 (_3I4489_$1I4488_$1I4620_SSRA, _3I4489_$1I4488_$1I4620_SSRA__vlIN);

 wire  _3I4489_$1I4488_$1I4620_SSRB;
 reg [1:16] _3I4489_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1206 (_3I4489_$1I4488_$1I4620_SSRB, _3I4489_$1I4488_$1I4620_SSRB__vlIN);

 wire  _3I4489_$1I4488_$1I4620_WEA;
 reg [1:16] _3I4489_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1207 (_3I4489_$1I4488_$1I4620_WEA, _3I4489_$1I4488_$1I4620_WEA__vlIN);

 wire  _3I4489_$1I4488_$1I4620_WEB;
 reg [1:16] _3I4489_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1208 (_3I4489_$1I4488_$1I4620_WEB, _3I4489_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _3I4489_$1I4488_$1I4620 ( _3I4489_$1I4488_$1I4620_DOA , _3I4489_$1I4488_$1I4620_DOB , _3I4489_$1I4488_$1I4620_DOPA , _3I4489_$1I4488_$1I4620_DOPB , _3I4489_$1I4488_$1I4620_ADDRA , _3I4489_$1I4488_$1I4620_ADDRB , _3I4489_$1I4488_$1I4620_CLKA , _3I4489_$1I4488_$1I4620_CLKB , _3I4489_$1I4488_$1I4620_DIA , _3I4489_$1I4488_$1I4620_DIB , _3I4489_$1I4488_$1I4620_DIPA , _3I4489_$1I4488_$1I4620_DIPB , _3I4489_$1I4488_$1I4620_ENA , _3I4489_$1I4488_$1I4620_ENB , _3I4489_$1I4488_$1I4620_SSRA , _3I4489_$1I4488_$1I4620_SSRB , _3I4489_$1I4488_$1I4620_WEA , _3I4489_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4464_$1I4488_$1I4621_DOA;

 wire [15:0] _3I4464_$1I4488_$1I4621_DOB;

 wire [0:0] _3I4464_$1I4488_$1I4621_DOPA;

 wire [1:0] _3I4464_$1I4488_$1I4621_DOPB;

 wire [10:0] _3I4464_$1I4488_$1I4621_ADDRA;
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1209_10 (_3I4464_$1I4488_$1I4621_ADDRA[10], _3I4464_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1209_9 (_3I4464_$1I4488_$1I4621_ADDRA[9], _3I4464_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1209_8 (_3I4464_$1I4488_$1I4621_ADDRA[8], _3I4464_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1209_7 (_3I4464_$1I4488_$1I4621_ADDRA[7], _3I4464_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1209_6 (_3I4464_$1I4488_$1I4621_ADDRA[6], _3I4464_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1209_5 (_3I4464_$1I4488_$1I4621_ADDRA[5], _3I4464_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1209_4 (_3I4464_$1I4488_$1I4621_ADDRA[4], _3I4464_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1209_3 (_3I4464_$1I4488_$1I4621_ADDRA[3], _3I4464_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1209_2 (_3I4464_$1I4488_$1I4621_ADDRA[2], _3I4464_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1209_1 (_3I4464_$1I4488_$1I4621_ADDRA[1], _3I4464_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1209_0 (_3I4464_$1I4488_$1I4621_ADDRA[0], _3I4464_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _3I4464_$1I4488_$1I4621_ADDRB;
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_1210_9 (_3I4464_$1I4488_$1I4621_ADDRB[9], _3I4464_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_1210_8 (_3I4464_$1I4488_$1I4621_ADDRB[8], _3I4464_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_1210_7 (_3I4464_$1I4488_$1I4621_ADDRB[7], _3I4464_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_1210_6 (_3I4464_$1I4488_$1I4621_ADDRB[6], _3I4464_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_1210_5 (_3I4464_$1I4488_$1I4621_ADDRB[5], _3I4464_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_1210_4 (_3I4464_$1I4488_$1I4621_ADDRB[4], _3I4464_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_1210_3 (_3I4464_$1I4488_$1I4621_ADDRB[3], _3I4464_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_1210_2 (_3I4464_$1I4488_$1I4621_ADDRB[2], _3I4464_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_1210_1 (_3I4464_$1I4488_$1I4621_ADDRB[1], _3I4464_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_1210_0 (_3I4464_$1I4488_$1I4621_ADDRB[0], _3I4464_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _3I4464_$1I4488_$1I4621_CLKA;
 reg [1:16] _3I4464_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_1211 (_3I4464_$1I4488_$1I4621_CLKA, _3I4464_$1I4488_$1I4621_CLKA__vlIN);

 wire  _3I4464_$1I4488_$1I4621_CLKB;
 reg [1:16] _3I4464_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_1212 (_3I4464_$1I4488_$1I4621_CLKB, _3I4464_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _3I4464_$1I4488_$1I4621_DIA;
 reg [1:16] _3I4464_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_1213_7 (_3I4464_$1I4488_$1I4621_DIA[7], _3I4464_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_1213_6 (_3I4464_$1I4488_$1I4621_DIA[6], _3I4464_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_1213_5 (_3I4464_$1I4488_$1I4621_DIA[5], _3I4464_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_1213_4 (_3I4464_$1I4488_$1I4621_DIA[4], _3I4464_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_1213_3 (_3I4464_$1I4488_$1I4621_DIA[3], _3I4464_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_1213_2 (_3I4464_$1I4488_$1I4621_DIA[2], _3I4464_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_1213_1 (_3I4464_$1I4488_$1I4621_DIA[1], _3I4464_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_1213_0 (_3I4464_$1I4488_$1I4621_DIA[0], _3I4464_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _3I4464_$1I4488_$1I4621_DIB;
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_1214_15 (_3I4464_$1I4488_$1I4621_DIB[15], _3I4464_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_1214_14 (_3I4464_$1I4488_$1I4621_DIB[14], _3I4464_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_1214_13 (_3I4464_$1I4488_$1I4621_DIB[13], _3I4464_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_1214_12 (_3I4464_$1I4488_$1I4621_DIB[12], _3I4464_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_1214_11 (_3I4464_$1I4488_$1I4621_DIB[11], _3I4464_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_1214_10 (_3I4464_$1I4488_$1I4621_DIB[10], _3I4464_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_1214_9 (_3I4464_$1I4488_$1I4621_DIB[9], _3I4464_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_1214_8 (_3I4464_$1I4488_$1I4621_DIB[8], _3I4464_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_1214_7 (_3I4464_$1I4488_$1I4621_DIB[7], _3I4464_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_1214_6 (_3I4464_$1I4488_$1I4621_DIB[6], _3I4464_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_1214_5 (_3I4464_$1I4488_$1I4621_DIB[5], _3I4464_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_1214_4 (_3I4464_$1I4488_$1I4621_DIB[4], _3I4464_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_1214_3 (_3I4464_$1I4488_$1I4621_DIB[3], _3I4464_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_1214_2 (_3I4464_$1I4488_$1I4621_DIB[2], _3I4464_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_1214_1 (_3I4464_$1I4488_$1I4621_DIB[1], _3I4464_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_1214_0 (_3I4464_$1I4488_$1I4621_DIB[0], _3I4464_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _3I4464_$1I4488_$1I4621_DIPA;
 reg [1:16] _3I4464_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_1215_0 (_3I4464_$1I4488_$1I4621_DIPA[0], _3I4464_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _3I4464_$1I4488_$1I4621_DIPB;
 reg [1:16] _3I4464_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_1216_1 (_3I4464_$1I4488_$1I4621_DIPB[1], _3I4464_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_1216_0 (_3I4464_$1I4488_$1I4621_DIPB[0], _3I4464_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _3I4464_$1I4488_$1I4621_ENA;
 reg [1:16] _3I4464_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_1217 (_3I4464_$1I4488_$1I4621_ENA, _3I4464_$1I4488_$1I4621_ENA__vlIN);

 wire  _3I4464_$1I4488_$1I4621_ENB;
 reg [1:16] _3I4464_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_1218 (_3I4464_$1I4488_$1I4621_ENB, _3I4464_$1I4488_$1I4621_ENB__vlIN);

 wire  _3I4464_$1I4488_$1I4621_SSRA;
 reg [1:16] _3I4464_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_1219 (_3I4464_$1I4488_$1I4621_SSRA, _3I4464_$1I4488_$1I4621_SSRA__vlIN);

 wire  _3I4464_$1I4488_$1I4621_SSRB;
 reg [1:16] _3I4464_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_1220 (_3I4464_$1I4488_$1I4621_SSRB, _3I4464_$1I4488_$1I4621_SSRB__vlIN);

 wire  _3I4464_$1I4488_$1I4621_WEA;
 reg [1:16] _3I4464_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_1221 (_3I4464_$1I4488_$1I4621_WEA, _3I4464_$1I4488_$1I4621_WEA__vlIN);

 wire  _3I4464_$1I4488_$1I4621_WEB;
 reg [1:16] _3I4464_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_1222 (_3I4464_$1I4488_$1I4621_WEB, _3I4464_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _3I4464_$1I4488_$1I4621 ( _3I4464_$1I4488_$1I4621_DOA , _3I4464_$1I4488_$1I4621_DOB , _3I4464_$1I4488_$1I4621_DOPA , _3I4464_$1I4488_$1I4621_DOPB , _3I4464_$1I4488_$1I4621_ADDRA , _3I4464_$1I4488_$1I4621_ADDRB , _3I4464_$1I4488_$1I4621_CLKA , _3I4464_$1I4488_$1I4621_CLKB , _3I4464_$1I4488_$1I4621_DIA , _3I4464_$1I4488_$1I4621_DIB , _3I4464_$1I4488_$1I4621_DIPA , _3I4464_$1I4488_$1I4621_DIPB , _3I4464_$1I4488_$1I4621_ENA , _3I4464_$1I4488_$1I4621_ENB , _3I4464_$1I4488_$1I4621_SSRA , _3I4464_$1I4488_$1I4621_SSRB , _3I4464_$1I4488_$1I4621_WEA , _3I4464_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4464_$1I4488_$1I4620_DOA;

 wire [15:0] _3I4464_$1I4488_$1I4620_DOB;

 wire [0:0] _3I4464_$1I4488_$1I4620_DOPA;

 wire [1:0] _3I4464_$1I4488_$1I4620_DOPB;

 wire [10:0] _3I4464_$1I4488_$1I4620_ADDRA;
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_1223_10 (_3I4464_$1I4488_$1I4620_ADDRA[10], _3I4464_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_1223_9 (_3I4464_$1I4488_$1I4620_ADDRA[9], _3I4464_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_1223_8 (_3I4464_$1I4488_$1I4620_ADDRA[8], _3I4464_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_1223_7 (_3I4464_$1I4488_$1I4620_ADDRA[7], _3I4464_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_1223_6 (_3I4464_$1I4488_$1I4620_ADDRA[6], _3I4464_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_1223_5 (_3I4464_$1I4488_$1I4620_ADDRA[5], _3I4464_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_1223_4 (_3I4464_$1I4488_$1I4620_ADDRA[4], _3I4464_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_1223_3 (_3I4464_$1I4488_$1I4620_ADDRA[3], _3I4464_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_1223_2 (_3I4464_$1I4488_$1I4620_ADDRA[2], _3I4464_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_1223_1 (_3I4464_$1I4488_$1I4620_ADDRA[1], _3I4464_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_1223_0 (_3I4464_$1I4488_$1I4620_ADDRA[0], _3I4464_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _3I4464_$1I4488_$1I4620_ADDRB;
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1224_9 (_3I4464_$1I4488_$1I4620_ADDRB[9], _3I4464_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1224_8 (_3I4464_$1I4488_$1I4620_ADDRB[8], _3I4464_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1224_7 (_3I4464_$1I4488_$1I4620_ADDRB[7], _3I4464_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1224_6 (_3I4464_$1I4488_$1I4620_ADDRB[6], _3I4464_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1224_5 (_3I4464_$1I4488_$1I4620_ADDRB[5], _3I4464_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1224_4 (_3I4464_$1I4488_$1I4620_ADDRB[4], _3I4464_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1224_3 (_3I4464_$1I4488_$1I4620_ADDRB[3], _3I4464_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1224_2 (_3I4464_$1I4488_$1I4620_ADDRB[2], _3I4464_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1224_1 (_3I4464_$1I4488_$1I4620_ADDRB[1], _3I4464_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1224_0 (_3I4464_$1I4488_$1I4620_ADDRB[0], _3I4464_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _3I4464_$1I4488_$1I4620_CLKA;
 reg [1:16] _3I4464_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1225 (_3I4464_$1I4488_$1I4620_CLKA, _3I4464_$1I4488_$1I4620_CLKA__vlIN);

 wire  _3I4464_$1I4488_$1I4620_CLKB;
 reg [1:16] _3I4464_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1226 (_3I4464_$1I4488_$1I4620_CLKB, _3I4464_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _3I4464_$1I4488_$1I4620_DIA;
 reg [1:16] _3I4464_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1227_7 (_3I4464_$1I4488_$1I4620_DIA[7], _3I4464_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1227_6 (_3I4464_$1I4488_$1I4620_DIA[6], _3I4464_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1227_5 (_3I4464_$1I4488_$1I4620_DIA[5], _3I4464_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1227_4 (_3I4464_$1I4488_$1I4620_DIA[4], _3I4464_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1227_3 (_3I4464_$1I4488_$1I4620_DIA[3], _3I4464_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1227_2 (_3I4464_$1I4488_$1I4620_DIA[2], _3I4464_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1227_1 (_3I4464_$1I4488_$1I4620_DIA[1], _3I4464_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1227_0 (_3I4464_$1I4488_$1I4620_DIA[0], _3I4464_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _3I4464_$1I4488_$1I4620_DIB;
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1228_15 (_3I4464_$1I4488_$1I4620_DIB[15], _3I4464_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1228_14 (_3I4464_$1I4488_$1I4620_DIB[14], _3I4464_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1228_13 (_3I4464_$1I4488_$1I4620_DIB[13], _3I4464_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1228_12 (_3I4464_$1I4488_$1I4620_DIB[12], _3I4464_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1228_11 (_3I4464_$1I4488_$1I4620_DIB[11], _3I4464_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1228_10 (_3I4464_$1I4488_$1I4620_DIB[10], _3I4464_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1228_9 (_3I4464_$1I4488_$1I4620_DIB[9], _3I4464_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1228_8 (_3I4464_$1I4488_$1I4620_DIB[8], _3I4464_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1228_7 (_3I4464_$1I4488_$1I4620_DIB[7], _3I4464_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1228_6 (_3I4464_$1I4488_$1I4620_DIB[6], _3I4464_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1228_5 (_3I4464_$1I4488_$1I4620_DIB[5], _3I4464_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1228_4 (_3I4464_$1I4488_$1I4620_DIB[4], _3I4464_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1228_3 (_3I4464_$1I4488_$1I4620_DIB[3], _3I4464_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1228_2 (_3I4464_$1I4488_$1I4620_DIB[2], _3I4464_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1228_1 (_3I4464_$1I4488_$1I4620_DIB[1], _3I4464_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1228_0 (_3I4464_$1I4488_$1I4620_DIB[0], _3I4464_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _3I4464_$1I4488_$1I4620_DIPA;
 reg [1:16] _3I4464_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1229_0 (_3I4464_$1I4488_$1I4620_DIPA[0], _3I4464_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _3I4464_$1I4488_$1I4620_DIPB;
 reg [1:16] _3I4464_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1230_1 (_3I4464_$1I4488_$1I4620_DIPB[1], _3I4464_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _3I4464_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1230_0 (_3I4464_$1I4488_$1I4620_DIPB[0], _3I4464_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _3I4464_$1I4488_$1I4620_ENA;
 reg [1:16] _3I4464_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1231 (_3I4464_$1I4488_$1I4620_ENA, _3I4464_$1I4488_$1I4620_ENA__vlIN);

 wire  _3I4464_$1I4488_$1I4620_ENB;
 reg [1:16] _3I4464_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1232 (_3I4464_$1I4488_$1I4620_ENB, _3I4464_$1I4488_$1I4620_ENB__vlIN);

 wire  _3I4464_$1I4488_$1I4620_SSRA;
 reg [1:16] _3I4464_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1233 (_3I4464_$1I4488_$1I4620_SSRA, _3I4464_$1I4488_$1I4620_SSRA__vlIN);

 wire  _3I4464_$1I4488_$1I4620_SSRB;
 reg [1:16] _3I4464_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1234 (_3I4464_$1I4488_$1I4620_SSRB, _3I4464_$1I4488_$1I4620_SSRB__vlIN);

 wire  _3I4464_$1I4488_$1I4620_WEA;
 reg [1:16] _3I4464_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1235 (_3I4464_$1I4488_$1I4620_WEA, _3I4464_$1I4488_$1I4620_WEA__vlIN);

 wire  _3I4464_$1I4488_$1I4620_WEB;
 reg [1:16] _3I4464_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1236 (_3I4464_$1I4488_$1I4620_WEB, _3I4464_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _3I4464_$1I4488_$1I4620 ( _3I4464_$1I4488_$1I4620_DOA , _3I4464_$1I4488_$1I4620_DOB , _3I4464_$1I4488_$1I4620_DOPA , _3I4464_$1I4488_$1I4620_DOPB , _3I4464_$1I4488_$1I4620_ADDRA , _3I4464_$1I4488_$1I4620_ADDRB , _3I4464_$1I4488_$1I4620_CLKA , _3I4464_$1I4488_$1I4620_CLKB , _3I4464_$1I4488_$1I4620_DIA , _3I4464_$1I4488_$1I4620_DIB , _3I4464_$1I4488_$1I4620_DIPA , _3I4464_$1I4488_$1I4620_DIPB , _3I4464_$1I4488_$1I4620_ENA , _3I4464_$1I4488_$1I4620_ENB , _3I4464_$1I4488_$1I4620_SSRA , _3I4464_$1I4488_$1I4620_SSRB , _3I4464_$1I4488_$1I4620_WEA , _3I4464_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4417_$1I4488_$1I4621_DOA;

 wire [15:0] _3I4417_$1I4488_$1I4621_DOB;

 wire [0:0] _3I4417_$1I4488_$1I4621_DOPA;

 wire [1:0] _3I4417_$1I4488_$1I4621_DOPB;

 wire [10:0] _3I4417_$1I4488_$1I4621_ADDRA;
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1237_10 (_3I4417_$1I4488_$1I4621_ADDRA[10], _3I4417_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1237_9 (_3I4417_$1I4488_$1I4621_ADDRA[9], _3I4417_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1237_8 (_3I4417_$1I4488_$1I4621_ADDRA[8], _3I4417_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1237_7 (_3I4417_$1I4488_$1I4621_ADDRA[7], _3I4417_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1237_6 (_3I4417_$1I4488_$1I4621_ADDRA[6], _3I4417_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1237_5 (_3I4417_$1I4488_$1I4621_ADDRA[5], _3I4417_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1237_4 (_3I4417_$1I4488_$1I4621_ADDRA[4], _3I4417_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1237_3 (_3I4417_$1I4488_$1I4621_ADDRA[3], _3I4417_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1237_2 (_3I4417_$1I4488_$1I4621_ADDRA[2], _3I4417_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1237_1 (_3I4417_$1I4488_$1I4621_ADDRA[1], _3I4417_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1237_0 (_3I4417_$1I4488_$1I4621_ADDRA[0], _3I4417_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _3I4417_$1I4488_$1I4621_ADDRB;
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_1238_9 (_3I4417_$1I4488_$1I4621_ADDRB[9], _3I4417_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_1238_8 (_3I4417_$1I4488_$1I4621_ADDRB[8], _3I4417_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_1238_7 (_3I4417_$1I4488_$1I4621_ADDRB[7], _3I4417_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_1238_6 (_3I4417_$1I4488_$1I4621_ADDRB[6], _3I4417_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_1238_5 (_3I4417_$1I4488_$1I4621_ADDRB[5], _3I4417_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_1238_4 (_3I4417_$1I4488_$1I4621_ADDRB[4], _3I4417_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_1238_3 (_3I4417_$1I4488_$1I4621_ADDRB[3], _3I4417_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_1238_2 (_3I4417_$1I4488_$1I4621_ADDRB[2], _3I4417_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_1238_1 (_3I4417_$1I4488_$1I4621_ADDRB[1], _3I4417_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_1238_0 (_3I4417_$1I4488_$1I4621_ADDRB[0], _3I4417_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _3I4417_$1I4488_$1I4621_CLKA;
 reg [1:16] _3I4417_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_1239 (_3I4417_$1I4488_$1I4621_CLKA, _3I4417_$1I4488_$1I4621_CLKA__vlIN);

 wire  _3I4417_$1I4488_$1I4621_CLKB;
 reg [1:16] _3I4417_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_1240 (_3I4417_$1I4488_$1I4621_CLKB, _3I4417_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _3I4417_$1I4488_$1I4621_DIA;
 reg [1:16] _3I4417_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_1241_7 (_3I4417_$1I4488_$1I4621_DIA[7], _3I4417_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_1241_6 (_3I4417_$1I4488_$1I4621_DIA[6], _3I4417_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_1241_5 (_3I4417_$1I4488_$1I4621_DIA[5], _3I4417_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_1241_4 (_3I4417_$1I4488_$1I4621_DIA[4], _3I4417_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_1241_3 (_3I4417_$1I4488_$1I4621_DIA[3], _3I4417_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_1241_2 (_3I4417_$1I4488_$1I4621_DIA[2], _3I4417_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_1241_1 (_3I4417_$1I4488_$1I4621_DIA[1], _3I4417_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_1241_0 (_3I4417_$1I4488_$1I4621_DIA[0], _3I4417_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _3I4417_$1I4488_$1I4621_DIB;
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_1242_15 (_3I4417_$1I4488_$1I4621_DIB[15], _3I4417_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_1242_14 (_3I4417_$1I4488_$1I4621_DIB[14], _3I4417_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_1242_13 (_3I4417_$1I4488_$1I4621_DIB[13], _3I4417_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_1242_12 (_3I4417_$1I4488_$1I4621_DIB[12], _3I4417_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_1242_11 (_3I4417_$1I4488_$1I4621_DIB[11], _3I4417_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_1242_10 (_3I4417_$1I4488_$1I4621_DIB[10], _3I4417_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_1242_9 (_3I4417_$1I4488_$1I4621_DIB[9], _3I4417_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_1242_8 (_3I4417_$1I4488_$1I4621_DIB[8], _3I4417_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_1242_7 (_3I4417_$1I4488_$1I4621_DIB[7], _3I4417_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_1242_6 (_3I4417_$1I4488_$1I4621_DIB[6], _3I4417_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_1242_5 (_3I4417_$1I4488_$1I4621_DIB[5], _3I4417_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_1242_4 (_3I4417_$1I4488_$1I4621_DIB[4], _3I4417_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_1242_3 (_3I4417_$1I4488_$1I4621_DIB[3], _3I4417_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_1242_2 (_3I4417_$1I4488_$1I4621_DIB[2], _3I4417_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_1242_1 (_3I4417_$1I4488_$1I4621_DIB[1], _3I4417_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_1242_0 (_3I4417_$1I4488_$1I4621_DIB[0], _3I4417_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _3I4417_$1I4488_$1I4621_DIPA;
 reg [1:16] _3I4417_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_1243_0 (_3I4417_$1I4488_$1I4621_DIPA[0], _3I4417_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _3I4417_$1I4488_$1I4621_DIPB;
 reg [1:16] _3I4417_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_1244_1 (_3I4417_$1I4488_$1I4621_DIPB[1], _3I4417_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_1244_0 (_3I4417_$1I4488_$1I4621_DIPB[0], _3I4417_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _3I4417_$1I4488_$1I4621_ENA;
 reg [1:16] _3I4417_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_1245 (_3I4417_$1I4488_$1I4621_ENA, _3I4417_$1I4488_$1I4621_ENA__vlIN);

 wire  _3I4417_$1I4488_$1I4621_ENB;
 reg [1:16] _3I4417_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_1246 (_3I4417_$1I4488_$1I4621_ENB, _3I4417_$1I4488_$1I4621_ENB__vlIN);

 wire  _3I4417_$1I4488_$1I4621_SSRA;
 reg [1:16] _3I4417_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_1247 (_3I4417_$1I4488_$1I4621_SSRA, _3I4417_$1I4488_$1I4621_SSRA__vlIN);

 wire  _3I4417_$1I4488_$1I4621_SSRB;
 reg [1:16] _3I4417_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_1248 (_3I4417_$1I4488_$1I4621_SSRB, _3I4417_$1I4488_$1I4621_SSRB__vlIN);

 wire  _3I4417_$1I4488_$1I4621_WEA;
 reg [1:16] _3I4417_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_1249 (_3I4417_$1I4488_$1I4621_WEA, _3I4417_$1I4488_$1I4621_WEA__vlIN);

 wire  _3I4417_$1I4488_$1I4621_WEB;
 reg [1:16] _3I4417_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_1250 (_3I4417_$1I4488_$1I4621_WEB, _3I4417_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _3I4417_$1I4488_$1I4621 ( _3I4417_$1I4488_$1I4621_DOA , _3I4417_$1I4488_$1I4621_DOB , _3I4417_$1I4488_$1I4621_DOPA , _3I4417_$1I4488_$1I4621_DOPB , _3I4417_$1I4488_$1I4621_ADDRA , _3I4417_$1I4488_$1I4621_ADDRB , _3I4417_$1I4488_$1I4621_CLKA , _3I4417_$1I4488_$1I4621_CLKB , _3I4417_$1I4488_$1I4621_DIA , _3I4417_$1I4488_$1I4621_DIB , _3I4417_$1I4488_$1I4621_DIPA , _3I4417_$1I4488_$1I4621_DIPB , _3I4417_$1I4488_$1I4621_ENA , _3I4417_$1I4488_$1I4621_ENB , _3I4417_$1I4488_$1I4621_SSRA , _3I4417_$1I4488_$1I4621_SSRB , _3I4417_$1I4488_$1I4621_WEA , _3I4417_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4417_$1I4488_$1I4620_DOA;

 wire [15:0] _3I4417_$1I4488_$1I4620_DOB;

 wire [0:0] _3I4417_$1I4488_$1I4620_DOPA;

 wire [1:0] _3I4417_$1I4488_$1I4620_DOPB;

 wire [10:0] _3I4417_$1I4488_$1I4620_ADDRA;
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_1251_10 (_3I4417_$1I4488_$1I4620_ADDRA[10], _3I4417_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_1251_9 (_3I4417_$1I4488_$1I4620_ADDRA[9], _3I4417_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_1251_8 (_3I4417_$1I4488_$1I4620_ADDRA[8], _3I4417_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_1251_7 (_3I4417_$1I4488_$1I4620_ADDRA[7], _3I4417_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_1251_6 (_3I4417_$1I4488_$1I4620_ADDRA[6], _3I4417_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_1251_5 (_3I4417_$1I4488_$1I4620_ADDRA[5], _3I4417_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_1251_4 (_3I4417_$1I4488_$1I4620_ADDRA[4], _3I4417_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_1251_3 (_3I4417_$1I4488_$1I4620_ADDRA[3], _3I4417_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_1251_2 (_3I4417_$1I4488_$1I4620_ADDRA[2], _3I4417_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_1251_1 (_3I4417_$1I4488_$1I4620_ADDRA[1], _3I4417_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_1251_0 (_3I4417_$1I4488_$1I4620_ADDRA[0], _3I4417_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _3I4417_$1I4488_$1I4620_ADDRB;
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1252_9 (_3I4417_$1I4488_$1I4620_ADDRB[9], _3I4417_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1252_8 (_3I4417_$1I4488_$1I4620_ADDRB[8], _3I4417_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1252_7 (_3I4417_$1I4488_$1I4620_ADDRB[7], _3I4417_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1252_6 (_3I4417_$1I4488_$1I4620_ADDRB[6], _3I4417_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1252_5 (_3I4417_$1I4488_$1I4620_ADDRB[5], _3I4417_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1252_4 (_3I4417_$1I4488_$1I4620_ADDRB[4], _3I4417_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1252_3 (_3I4417_$1I4488_$1I4620_ADDRB[3], _3I4417_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1252_2 (_3I4417_$1I4488_$1I4620_ADDRB[2], _3I4417_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1252_1 (_3I4417_$1I4488_$1I4620_ADDRB[1], _3I4417_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1252_0 (_3I4417_$1I4488_$1I4620_ADDRB[0], _3I4417_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _3I4417_$1I4488_$1I4620_CLKA;
 reg [1:16] _3I4417_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1253 (_3I4417_$1I4488_$1I4620_CLKA, _3I4417_$1I4488_$1I4620_CLKA__vlIN);

 wire  _3I4417_$1I4488_$1I4620_CLKB;
 reg [1:16] _3I4417_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1254 (_3I4417_$1I4488_$1I4620_CLKB, _3I4417_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _3I4417_$1I4488_$1I4620_DIA;
 reg [1:16] _3I4417_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1255_7 (_3I4417_$1I4488_$1I4620_DIA[7], _3I4417_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1255_6 (_3I4417_$1I4488_$1I4620_DIA[6], _3I4417_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1255_5 (_3I4417_$1I4488_$1I4620_DIA[5], _3I4417_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1255_4 (_3I4417_$1I4488_$1I4620_DIA[4], _3I4417_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1255_3 (_3I4417_$1I4488_$1I4620_DIA[3], _3I4417_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1255_2 (_3I4417_$1I4488_$1I4620_DIA[2], _3I4417_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1255_1 (_3I4417_$1I4488_$1I4620_DIA[1], _3I4417_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1255_0 (_3I4417_$1I4488_$1I4620_DIA[0], _3I4417_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _3I4417_$1I4488_$1I4620_DIB;
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1256_15 (_3I4417_$1I4488_$1I4620_DIB[15], _3I4417_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1256_14 (_3I4417_$1I4488_$1I4620_DIB[14], _3I4417_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1256_13 (_3I4417_$1I4488_$1I4620_DIB[13], _3I4417_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1256_12 (_3I4417_$1I4488_$1I4620_DIB[12], _3I4417_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1256_11 (_3I4417_$1I4488_$1I4620_DIB[11], _3I4417_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1256_10 (_3I4417_$1I4488_$1I4620_DIB[10], _3I4417_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1256_9 (_3I4417_$1I4488_$1I4620_DIB[9], _3I4417_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1256_8 (_3I4417_$1I4488_$1I4620_DIB[8], _3I4417_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1256_7 (_3I4417_$1I4488_$1I4620_DIB[7], _3I4417_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1256_6 (_3I4417_$1I4488_$1I4620_DIB[6], _3I4417_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1256_5 (_3I4417_$1I4488_$1I4620_DIB[5], _3I4417_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1256_4 (_3I4417_$1I4488_$1I4620_DIB[4], _3I4417_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1256_3 (_3I4417_$1I4488_$1I4620_DIB[3], _3I4417_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1256_2 (_3I4417_$1I4488_$1I4620_DIB[2], _3I4417_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1256_1 (_3I4417_$1I4488_$1I4620_DIB[1], _3I4417_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1256_0 (_3I4417_$1I4488_$1I4620_DIB[0], _3I4417_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _3I4417_$1I4488_$1I4620_DIPA;
 reg [1:16] _3I4417_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1257_0 (_3I4417_$1I4488_$1I4620_DIPA[0], _3I4417_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _3I4417_$1I4488_$1I4620_DIPB;
 reg [1:16] _3I4417_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1258_1 (_3I4417_$1I4488_$1I4620_DIPB[1], _3I4417_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _3I4417_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1258_0 (_3I4417_$1I4488_$1I4620_DIPB[0], _3I4417_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _3I4417_$1I4488_$1I4620_ENA;
 reg [1:16] _3I4417_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1259 (_3I4417_$1I4488_$1I4620_ENA, _3I4417_$1I4488_$1I4620_ENA__vlIN);

 wire  _3I4417_$1I4488_$1I4620_ENB;
 reg [1:16] _3I4417_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1260 (_3I4417_$1I4488_$1I4620_ENB, _3I4417_$1I4488_$1I4620_ENB__vlIN);

 wire  _3I4417_$1I4488_$1I4620_SSRA;
 reg [1:16] _3I4417_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1261 (_3I4417_$1I4488_$1I4620_SSRA, _3I4417_$1I4488_$1I4620_SSRA__vlIN);

 wire  _3I4417_$1I4488_$1I4620_SSRB;
 reg [1:16] _3I4417_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1262 (_3I4417_$1I4488_$1I4620_SSRB, _3I4417_$1I4488_$1I4620_SSRB__vlIN);

 wire  _3I4417_$1I4488_$1I4620_WEA;
 reg [1:16] _3I4417_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1263 (_3I4417_$1I4488_$1I4620_WEA, _3I4417_$1I4488_$1I4620_WEA__vlIN);

 wire  _3I4417_$1I4488_$1I4620_WEB;
 reg [1:16] _3I4417_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1264 (_3I4417_$1I4488_$1I4620_WEB, _3I4417_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _3I4417_$1I4488_$1I4620 ( _3I4417_$1I4488_$1I4620_DOA , _3I4417_$1I4488_$1I4620_DOB , _3I4417_$1I4488_$1I4620_DOPA , _3I4417_$1I4488_$1I4620_DOPB , _3I4417_$1I4488_$1I4620_ADDRA , _3I4417_$1I4488_$1I4620_ADDRB , _3I4417_$1I4488_$1I4620_CLKA , _3I4417_$1I4488_$1I4620_CLKB , _3I4417_$1I4488_$1I4620_DIA , _3I4417_$1I4488_$1I4620_DIB , _3I4417_$1I4488_$1I4620_DIPA , _3I4417_$1I4488_$1I4620_DIPB , _3I4417_$1I4488_$1I4620_ENA , _3I4417_$1I4488_$1I4620_ENB , _3I4417_$1I4488_$1I4620_SSRA , _3I4417_$1I4488_$1I4620_SSRB , _3I4417_$1I4488_$1I4620_WEA , _3I4417_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4392_$1I4488_$1I4621_DOA;

 wire [15:0] _3I4392_$1I4488_$1I4621_DOB;

 wire [0:0] _3I4392_$1I4488_$1I4621_DOPA;

 wire [1:0] _3I4392_$1I4488_$1I4621_DOPB;

 wire [10:0] _3I4392_$1I4488_$1I4621_ADDRA;
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1265_10 (_3I4392_$1I4488_$1I4621_ADDRA[10], _3I4392_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1265_9 (_3I4392_$1I4488_$1I4621_ADDRA[9], _3I4392_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1265_8 (_3I4392_$1I4488_$1I4621_ADDRA[8], _3I4392_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1265_7 (_3I4392_$1I4488_$1I4621_ADDRA[7], _3I4392_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1265_6 (_3I4392_$1I4488_$1I4621_ADDRA[6], _3I4392_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1265_5 (_3I4392_$1I4488_$1I4621_ADDRA[5], _3I4392_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1265_4 (_3I4392_$1I4488_$1I4621_ADDRA[4], _3I4392_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1265_3 (_3I4392_$1I4488_$1I4621_ADDRA[3], _3I4392_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1265_2 (_3I4392_$1I4488_$1I4621_ADDRA[2], _3I4392_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1265_1 (_3I4392_$1I4488_$1I4621_ADDRA[1], _3I4392_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1265_0 (_3I4392_$1I4488_$1I4621_ADDRA[0], _3I4392_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _3I4392_$1I4488_$1I4621_ADDRB;
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_1266_9 (_3I4392_$1I4488_$1I4621_ADDRB[9], _3I4392_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_1266_8 (_3I4392_$1I4488_$1I4621_ADDRB[8], _3I4392_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_1266_7 (_3I4392_$1I4488_$1I4621_ADDRB[7], _3I4392_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_1266_6 (_3I4392_$1I4488_$1I4621_ADDRB[6], _3I4392_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_1266_5 (_3I4392_$1I4488_$1I4621_ADDRB[5], _3I4392_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_1266_4 (_3I4392_$1I4488_$1I4621_ADDRB[4], _3I4392_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_1266_3 (_3I4392_$1I4488_$1I4621_ADDRB[3], _3I4392_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_1266_2 (_3I4392_$1I4488_$1I4621_ADDRB[2], _3I4392_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_1266_1 (_3I4392_$1I4488_$1I4621_ADDRB[1], _3I4392_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_1266_0 (_3I4392_$1I4488_$1I4621_ADDRB[0], _3I4392_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _3I4392_$1I4488_$1I4621_CLKA;
 reg [1:16] _3I4392_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_1267 (_3I4392_$1I4488_$1I4621_CLKA, _3I4392_$1I4488_$1I4621_CLKA__vlIN);

 wire  _3I4392_$1I4488_$1I4621_CLKB;
 reg [1:16] _3I4392_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_1268 (_3I4392_$1I4488_$1I4621_CLKB, _3I4392_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _3I4392_$1I4488_$1I4621_DIA;
 reg [1:16] _3I4392_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_1269_7 (_3I4392_$1I4488_$1I4621_DIA[7], _3I4392_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_1269_6 (_3I4392_$1I4488_$1I4621_DIA[6], _3I4392_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_1269_5 (_3I4392_$1I4488_$1I4621_DIA[5], _3I4392_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_1269_4 (_3I4392_$1I4488_$1I4621_DIA[4], _3I4392_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_1269_3 (_3I4392_$1I4488_$1I4621_DIA[3], _3I4392_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_1269_2 (_3I4392_$1I4488_$1I4621_DIA[2], _3I4392_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_1269_1 (_3I4392_$1I4488_$1I4621_DIA[1], _3I4392_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_1269_0 (_3I4392_$1I4488_$1I4621_DIA[0], _3I4392_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _3I4392_$1I4488_$1I4621_DIB;
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_1270_15 (_3I4392_$1I4488_$1I4621_DIB[15], _3I4392_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_1270_14 (_3I4392_$1I4488_$1I4621_DIB[14], _3I4392_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_1270_13 (_3I4392_$1I4488_$1I4621_DIB[13], _3I4392_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_1270_12 (_3I4392_$1I4488_$1I4621_DIB[12], _3I4392_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_1270_11 (_3I4392_$1I4488_$1I4621_DIB[11], _3I4392_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_1270_10 (_3I4392_$1I4488_$1I4621_DIB[10], _3I4392_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_1270_9 (_3I4392_$1I4488_$1I4621_DIB[9], _3I4392_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_1270_8 (_3I4392_$1I4488_$1I4621_DIB[8], _3I4392_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_1270_7 (_3I4392_$1I4488_$1I4621_DIB[7], _3I4392_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_1270_6 (_3I4392_$1I4488_$1I4621_DIB[6], _3I4392_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_1270_5 (_3I4392_$1I4488_$1I4621_DIB[5], _3I4392_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_1270_4 (_3I4392_$1I4488_$1I4621_DIB[4], _3I4392_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_1270_3 (_3I4392_$1I4488_$1I4621_DIB[3], _3I4392_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_1270_2 (_3I4392_$1I4488_$1I4621_DIB[2], _3I4392_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_1270_1 (_3I4392_$1I4488_$1I4621_DIB[1], _3I4392_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_1270_0 (_3I4392_$1I4488_$1I4621_DIB[0], _3I4392_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _3I4392_$1I4488_$1I4621_DIPA;
 reg [1:16] _3I4392_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_1271_0 (_3I4392_$1I4488_$1I4621_DIPA[0], _3I4392_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _3I4392_$1I4488_$1I4621_DIPB;
 reg [1:16] _3I4392_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_1272_1 (_3I4392_$1I4488_$1I4621_DIPB[1], _3I4392_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_1272_0 (_3I4392_$1I4488_$1I4621_DIPB[0], _3I4392_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _3I4392_$1I4488_$1I4621_ENA;
 reg [1:16] _3I4392_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_1273 (_3I4392_$1I4488_$1I4621_ENA, _3I4392_$1I4488_$1I4621_ENA__vlIN);

 wire  _3I4392_$1I4488_$1I4621_ENB;
 reg [1:16] _3I4392_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_1274 (_3I4392_$1I4488_$1I4621_ENB, _3I4392_$1I4488_$1I4621_ENB__vlIN);

 wire  _3I4392_$1I4488_$1I4621_SSRA;
 reg [1:16] _3I4392_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_1275 (_3I4392_$1I4488_$1I4621_SSRA, _3I4392_$1I4488_$1I4621_SSRA__vlIN);

 wire  _3I4392_$1I4488_$1I4621_SSRB;
 reg [1:16] _3I4392_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_1276 (_3I4392_$1I4488_$1I4621_SSRB, _3I4392_$1I4488_$1I4621_SSRB__vlIN);

 wire  _3I4392_$1I4488_$1I4621_WEA;
 reg [1:16] _3I4392_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_1277 (_3I4392_$1I4488_$1I4621_WEA, _3I4392_$1I4488_$1I4621_WEA__vlIN);

 wire  _3I4392_$1I4488_$1I4621_WEB;
 reg [1:16] _3I4392_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_1278 (_3I4392_$1I4488_$1I4621_WEB, _3I4392_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _3I4392_$1I4488_$1I4621 ( _3I4392_$1I4488_$1I4621_DOA , _3I4392_$1I4488_$1I4621_DOB , _3I4392_$1I4488_$1I4621_DOPA , _3I4392_$1I4488_$1I4621_DOPB , _3I4392_$1I4488_$1I4621_ADDRA , _3I4392_$1I4488_$1I4621_ADDRB , _3I4392_$1I4488_$1I4621_CLKA , _3I4392_$1I4488_$1I4621_CLKB , _3I4392_$1I4488_$1I4621_DIA , _3I4392_$1I4488_$1I4621_DIB , _3I4392_$1I4488_$1I4621_DIPA , _3I4392_$1I4488_$1I4621_DIPB , _3I4392_$1I4488_$1I4621_ENA , _3I4392_$1I4488_$1I4621_ENB , _3I4392_$1I4488_$1I4621_SSRA , _3I4392_$1I4488_$1I4621_SSRB , _3I4392_$1I4488_$1I4621_WEA , _3I4392_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4392_$1I4488_$1I4620_DOA;

 wire [15:0] _3I4392_$1I4488_$1I4620_DOB;

 wire [0:0] _3I4392_$1I4488_$1I4620_DOPA;

 wire [1:0] _3I4392_$1I4488_$1I4620_DOPB;

 wire [10:0] _3I4392_$1I4488_$1I4620_ADDRA;
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_1279_10 (_3I4392_$1I4488_$1I4620_ADDRA[10], _3I4392_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_1279_9 (_3I4392_$1I4488_$1I4620_ADDRA[9], _3I4392_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_1279_8 (_3I4392_$1I4488_$1I4620_ADDRA[8], _3I4392_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_1279_7 (_3I4392_$1I4488_$1I4620_ADDRA[7], _3I4392_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_1279_6 (_3I4392_$1I4488_$1I4620_ADDRA[6], _3I4392_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_1279_5 (_3I4392_$1I4488_$1I4620_ADDRA[5], _3I4392_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_1279_4 (_3I4392_$1I4488_$1I4620_ADDRA[4], _3I4392_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_1279_3 (_3I4392_$1I4488_$1I4620_ADDRA[3], _3I4392_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_1279_2 (_3I4392_$1I4488_$1I4620_ADDRA[2], _3I4392_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_1279_1 (_3I4392_$1I4488_$1I4620_ADDRA[1], _3I4392_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_1279_0 (_3I4392_$1I4488_$1I4620_ADDRA[0], _3I4392_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _3I4392_$1I4488_$1I4620_ADDRB;
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1280_9 (_3I4392_$1I4488_$1I4620_ADDRB[9], _3I4392_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1280_8 (_3I4392_$1I4488_$1I4620_ADDRB[8], _3I4392_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1280_7 (_3I4392_$1I4488_$1I4620_ADDRB[7], _3I4392_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1280_6 (_3I4392_$1I4488_$1I4620_ADDRB[6], _3I4392_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1280_5 (_3I4392_$1I4488_$1I4620_ADDRB[5], _3I4392_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1280_4 (_3I4392_$1I4488_$1I4620_ADDRB[4], _3I4392_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1280_3 (_3I4392_$1I4488_$1I4620_ADDRB[3], _3I4392_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1280_2 (_3I4392_$1I4488_$1I4620_ADDRB[2], _3I4392_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1280_1 (_3I4392_$1I4488_$1I4620_ADDRB[1], _3I4392_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1280_0 (_3I4392_$1I4488_$1I4620_ADDRB[0], _3I4392_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _3I4392_$1I4488_$1I4620_CLKA;
 reg [1:16] _3I4392_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1281 (_3I4392_$1I4488_$1I4620_CLKA, _3I4392_$1I4488_$1I4620_CLKA__vlIN);

 wire  _3I4392_$1I4488_$1I4620_CLKB;
 reg [1:16] _3I4392_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1282 (_3I4392_$1I4488_$1I4620_CLKB, _3I4392_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _3I4392_$1I4488_$1I4620_DIA;
 reg [1:16] _3I4392_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1283_7 (_3I4392_$1I4488_$1I4620_DIA[7], _3I4392_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1283_6 (_3I4392_$1I4488_$1I4620_DIA[6], _3I4392_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1283_5 (_3I4392_$1I4488_$1I4620_DIA[5], _3I4392_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1283_4 (_3I4392_$1I4488_$1I4620_DIA[4], _3I4392_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1283_3 (_3I4392_$1I4488_$1I4620_DIA[3], _3I4392_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1283_2 (_3I4392_$1I4488_$1I4620_DIA[2], _3I4392_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1283_1 (_3I4392_$1I4488_$1I4620_DIA[1], _3I4392_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1283_0 (_3I4392_$1I4488_$1I4620_DIA[0], _3I4392_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _3I4392_$1I4488_$1I4620_DIB;
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1284_15 (_3I4392_$1I4488_$1I4620_DIB[15], _3I4392_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1284_14 (_3I4392_$1I4488_$1I4620_DIB[14], _3I4392_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1284_13 (_3I4392_$1I4488_$1I4620_DIB[13], _3I4392_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1284_12 (_3I4392_$1I4488_$1I4620_DIB[12], _3I4392_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1284_11 (_3I4392_$1I4488_$1I4620_DIB[11], _3I4392_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1284_10 (_3I4392_$1I4488_$1I4620_DIB[10], _3I4392_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1284_9 (_3I4392_$1I4488_$1I4620_DIB[9], _3I4392_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1284_8 (_3I4392_$1I4488_$1I4620_DIB[8], _3I4392_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1284_7 (_3I4392_$1I4488_$1I4620_DIB[7], _3I4392_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1284_6 (_3I4392_$1I4488_$1I4620_DIB[6], _3I4392_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1284_5 (_3I4392_$1I4488_$1I4620_DIB[5], _3I4392_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1284_4 (_3I4392_$1I4488_$1I4620_DIB[4], _3I4392_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1284_3 (_3I4392_$1I4488_$1I4620_DIB[3], _3I4392_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1284_2 (_3I4392_$1I4488_$1I4620_DIB[2], _3I4392_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1284_1 (_3I4392_$1I4488_$1I4620_DIB[1], _3I4392_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1284_0 (_3I4392_$1I4488_$1I4620_DIB[0], _3I4392_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _3I4392_$1I4488_$1I4620_DIPA;
 reg [1:16] _3I4392_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1285_0 (_3I4392_$1I4488_$1I4620_DIPA[0], _3I4392_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _3I4392_$1I4488_$1I4620_DIPB;
 reg [1:16] _3I4392_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1286_1 (_3I4392_$1I4488_$1I4620_DIPB[1], _3I4392_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _3I4392_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1286_0 (_3I4392_$1I4488_$1I4620_DIPB[0], _3I4392_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _3I4392_$1I4488_$1I4620_ENA;
 reg [1:16] _3I4392_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1287 (_3I4392_$1I4488_$1I4620_ENA, _3I4392_$1I4488_$1I4620_ENA__vlIN);

 wire  _3I4392_$1I4488_$1I4620_ENB;
 reg [1:16] _3I4392_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1288 (_3I4392_$1I4488_$1I4620_ENB, _3I4392_$1I4488_$1I4620_ENB__vlIN);

 wire  _3I4392_$1I4488_$1I4620_SSRA;
 reg [1:16] _3I4392_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1289 (_3I4392_$1I4488_$1I4620_SSRA, _3I4392_$1I4488_$1I4620_SSRA__vlIN);

 wire  _3I4392_$1I4488_$1I4620_SSRB;
 reg [1:16] _3I4392_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1290 (_3I4392_$1I4488_$1I4620_SSRB, _3I4392_$1I4488_$1I4620_SSRB__vlIN);

 wire  _3I4392_$1I4488_$1I4620_WEA;
 reg [1:16] _3I4392_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1291 (_3I4392_$1I4488_$1I4620_WEA, _3I4392_$1I4488_$1I4620_WEA__vlIN);

 wire  _3I4392_$1I4488_$1I4620_WEB;
 reg [1:16] _3I4392_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1292 (_3I4392_$1I4488_$1I4620_WEB, _3I4392_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _3I4392_$1I4488_$1I4620 ( _3I4392_$1I4488_$1I4620_DOA , _3I4392_$1I4488_$1I4620_DOB , _3I4392_$1I4488_$1I4620_DOPA , _3I4392_$1I4488_$1I4620_DOPB , _3I4392_$1I4488_$1I4620_ADDRA , _3I4392_$1I4488_$1I4620_ADDRB , _3I4392_$1I4488_$1I4620_CLKA , _3I4392_$1I4488_$1I4620_CLKB , _3I4392_$1I4488_$1I4620_DIA , _3I4392_$1I4488_$1I4620_DIB , _3I4392_$1I4488_$1I4620_DIPA , _3I4392_$1I4488_$1I4620_DIPB , _3I4392_$1I4488_$1I4620_ENA , _3I4392_$1I4488_$1I4620_ENB , _3I4392_$1I4488_$1I4620_SSRA , _3I4392_$1I4488_$1I4620_SSRB , _3I4392_$1I4488_$1I4620_WEA , _3I4392_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4365_$1I4488_$1I4621_DOA;

 wire [15:0] _3I4365_$1I4488_$1I4621_DOB;

 wire [0:0] _3I4365_$1I4488_$1I4621_DOPA;

 wire [1:0] _3I4365_$1I4488_$1I4621_DOPB;

 wire [10:0] _3I4365_$1I4488_$1I4621_ADDRA;
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1293_10 (_3I4365_$1I4488_$1I4621_ADDRA[10], _3I4365_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1293_9 (_3I4365_$1I4488_$1I4621_ADDRA[9], _3I4365_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1293_8 (_3I4365_$1I4488_$1I4621_ADDRA[8], _3I4365_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1293_7 (_3I4365_$1I4488_$1I4621_ADDRA[7], _3I4365_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1293_6 (_3I4365_$1I4488_$1I4621_ADDRA[6], _3I4365_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1293_5 (_3I4365_$1I4488_$1I4621_ADDRA[5], _3I4365_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1293_4 (_3I4365_$1I4488_$1I4621_ADDRA[4], _3I4365_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1293_3 (_3I4365_$1I4488_$1I4621_ADDRA[3], _3I4365_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1293_2 (_3I4365_$1I4488_$1I4621_ADDRA[2], _3I4365_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1293_1 (_3I4365_$1I4488_$1I4621_ADDRA[1], _3I4365_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1293_0 (_3I4365_$1I4488_$1I4621_ADDRA[0], _3I4365_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _3I4365_$1I4488_$1I4621_ADDRB;
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_1294_9 (_3I4365_$1I4488_$1I4621_ADDRB[9], _3I4365_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_1294_8 (_3I4365_$1I4488_$1I4621_ADDRB[8], _3I4365_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_1294_7 (_3I4365_$1I4488_$1I4621_ADDRB[7], _3I4365_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_1294_6 (_3I4365_$1I4488_$1I4621_ADDRB[6], _3I4365_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_1294_5 (_3I4365_$1I4488_$1I4621_ADDRB[5], _3I4365_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_1294_4 (_3I4365_$1I4488_$1I4621_ADDRB[4], _3I4365_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_1294_3 (_3I4365_$1I4488_$1I4621_ADDRB[3], _3I4365_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_1294_2 (_3I4365_$1I4488_$1I4621_ADDRB[2], _3I4365_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_1294_1 (_3I4365_$1I4488_$1I4621_ADDRB[1], _3I4365_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_1294_0 (_3I4365_$1I4488_$1I4621_ADDRB[0], _3I4365_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _3I4365_$1I4488_$1I4621_CLKA;
 reg [1:16] _3I4365_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_1295 (_3I4365_$1I4488_$1I4621_CLKA, _3I4365_$1I4488_$1I4621_CLKA__vlIN);

 wire  _3I4365_$1I4488_$1I4621_CLKB;
 reg [1:16] _3I4365_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_1296 (_3I4365_$1I4488_$1I4621_CLKB, _3I4365_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _3I4365_$1I4488_$1I4621_DIA;
 reg [1:16] _3I4365_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_1297_7 (_3I4365_$1I4488_$1I4621_DIA[7], _3I4365_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_1297_6 (_3I4365_$1I4488_$1I4621_DIA[6], _3I4365_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_1297_5 (_3I4365_$1I4488_$1I4621_DIA[5], _3I4365_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_1297_4 (_3I4365_$1I4488_$1I4621_DIA[4], _3I4365_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_1297_3 (_3I4365_$1I4488_$1I4621_DIA[3], _3I4365_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_1297_2 (_3I4365_$1I4488_$1I4621_DIA[2], _3I4365_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_1297_1 (_3I4365_$1I4488_$1I4621_DIA[1], _3I4365_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_1297_0 (_3I4365_$1I4488_$1I4621_DIA[0], _3I4365_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _3I4365_$1I4488_$1I4621_DIB;
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_1298_15 (_3I4365_$1I4488_$1I4621_DIB[15], _3I4365_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_1298_14 (_3I4365_$1I4488_$1I4621_DIB[14], _3I4365_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_1298_13 (_3I4365_$1I4488_$1I4621_DIB[13], _3I4365_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_1298_12 (_3I4365_$1I4488_$1I4621_DIB[12], _3I4365_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_1298_11 (_3I4365_$1I4488_$1I4621_DIB[11], _3I4365_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_1298_10 (_3I4365_$1I4488_$1I4621_DIB[10], _3I4365_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_1298_9 (_3I4365_$1I4488_$1I4621_DIB[9], _3I4365_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_1298_8 (_3I4365_$1I4488_$1I4621_DIB[8], _3I4365_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_1298_7 (_3I4365_$1I4488_$1I4621_DIB[7], _3I4365_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_1298_6 (_3I4365_$1I4488_$1I4621_DIB[6], _3I4365_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_1298_5 (_3I4365_$1I4488_$1I4621_DIB[5], _3I4365_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_1298_4 (_3I4365_$1I4488_$1I4621_DIB[4], _3I4365_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_1298_3 (_3I4365_$1I4488_$1I4621_DIB[3], _3I4365_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_1298_2 (_3I4365_$1I4488_$1I4621_DIB[2], _3I4365_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_1298_1 (_3I4365_$1I4488_$1I4621_DIB[1], _3I4365_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_1298_0 (_3I4365_$1I4488_$1I4621_DIB[0], _3I4365_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _3I4365_$1I4488_$1I4621_DIPA;
 reg [1:16] _3I4365_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_1299_0 (_3I4365_$1I4488_$1I4621_DIPA[0], _3I4365_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _3I4365_$1I4488_$1I4621_DIPB;
 reg [1:16] _3I4365_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_1300_1 (_3I4365_$1I4488_$1I4621_DIPB[1], _3I4365_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_1300_0 (_3I4365_$1I4488_$1I4621_DIPB[0], _3I4365_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _3I4365_$1I4488_$1I4621_ENA;
 reg [1:16] _3I4365_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_1301 (_3I4365_$1I4488_$1I4621_ENA, _3I4365_$1I4488_$1I4621_ENA__vlIN);

 wire  _3I4365_$1I4488_$1I4621_ENB;
 reg [1:16] _3I4365_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_1302 (_3I4365_$1I4488_$1I4621_ENB, _3I4365_$1I4488_$1I4621_ENB__vlIN);

 wire  _3I4365_$1I4488_$1I4621_SSRA;
 reg [1:16] _3I4365_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_1303 (_3I4365_$1I4488_$1I4621_SSRA, _3I4365_$1I4488_$1I4621_SSRA__vlIN);

 wire  _3I4365_$1I4488_$1I4621_SSRB;
 reg [1:16] _3I4365_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_1304 (_3I4365_$1I4488_$1I4621_SSRB, _3I4365_$1I4488_$1I4621_SSRB__vlIN);

 wire  _3I4365_$1I4488_$1I4621_WEA;
 reg [1:16] _3I4365_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_1305 (_3I4365_$1I4488_$1I4621_WEA, _3I4365_$1I4488_$1I4621_WEA__vlIN);

 wire  _3I4365_$1I4488_$1I4621_WEB;
 reg [1:16] _3I4365_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_1306 (_3I4365_$1I4488_$1I4621_WEB, _3I4365_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _3I4365_$1I4488_$1I4621 ( _3I4365_$1I4488_$1I4621_DOA , _3I4365_$1I4488_$1I4621_DOB , _3I4365_$1I4488_$1I4621_DOPA , _3I4365_$1I4488_$1I4621_DOPB , _3I4365_$1I4488_$1I4621_ADDRA , _3I4365_$1I4488_$1I4621_ADDRB , _3I4365_$1I4488_$1I4621_CLKA , _3I4365_$1I4488_$1I4621_CLKB , _3I4365_$1I4488_$1I4621_DIA , _3I4365_$1I4488_$1I4621_DIB , _3I4365_$1I4488_$1I4621_DIPA , _3I4365_$1I4488_$1I4621_DIPB , _3I4365_$1I4488_$1I4621_ENA , _3I4365_$1I4488_$1I4621_ENB , _3I4365_$1I4488_$1I4621_SSRA , _3I4365_$1I4488_$1I4621_SSRB , _3I4365_$1I4488_$1I4621_WEA , _3I4365_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4365_$1I4488_$1I4620_DOA;

 wire [15:0] _3I4365_$1I4488_$1I4620_DOB;

 wire [0:0] _3I4365_$1I4488_$1I4620_DOPA;

 wire [1:0] _3I4365_$1I4488_$1I4620_DOPB;

 wire [10:0] _3I4365_$1I4488_$1I4620_ADDRA;
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_1307_10 (_3I4365_$1I4488_$1I4620_ADDRA[10], _3I4365_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_1307_9 (_3I4365_$1I4488_$1I4620_ADDRA[9], _3I4365_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_1307_8 (_3I4365_$1I4488_$1I4620_ADDRA[8], _3I4365_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_1307_7 (_3I4365_$1I4488_$1I4620_ADDRA[7], _3I4365_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_1307_6 (_3I4365_$1I4488_$1I4620_ADDRA[6], _3I4365_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_1307_5 (_3I4365_$1I4488_$1I4620_ADDRA[5], _3I4365_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_1307_4 (_3I4365_$1I4488_$1I4620_ADDRA[4], _3I4365_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_1307_3 (_3I4365_$1I4488_$1I4620_ADDRA[3], _3I4365_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_1307_2 (_3I4365_$1I4488_$1I4620_ADDRA[2], _3I4365_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_1307_1 (_3I4365_$1I4488_$1I4620_ADDRA[1], _3I4365_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_1307_0 (_3I4365_$1I4488_$1I4620_ADDRA[0], _3I4365_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _3I4365_$1I4488_$1I4620_ADDRB;
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1308_9 (_3I4365_$1I4488_$1I4620_ADDRB[9], _3I4365_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1308_8 (_3I4365_$1I4488_$1I4620_ADDRB[8], _3I4365_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1308_7 (_3I4365_$1I4488_$1I4620_ADDRB[7], _3I4365_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1308_6 (_3I4365_$1I4488_$1I4620_ADDRB[6], _3I4365_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1308_5 (_3I4365_$1I4488_$1I4620_ADDRB[5], _3I4365_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1308_4 (_3I4365_$1I4488_$1I4620_ADDRB[4], _3I4365_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1308_3 (_3I4365_$1I4488_$1I4620_ADDRB[3], _3I4365_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1308_2 (_3I4365_$1I4488_$1I4620_ADDRB[2], _3I4365_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1308_1 (_3I4365_$1I4488_$1I4620_ADDRB[1], _3I4365_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1308_0 (_3I4365_$1I4488_$1I4620_ADDRB[0], _3I4365_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _3I4365_$1I4488_$1I4620_CLKA;
 reg [1:16] _3I4365_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1309 (_3I4365_$1I4488_$1I4620_CLKA, _3I4365_$1I4488_$1I4620_CLKA__vlIN);

 wire  _3I4365_$1I4488_$1I4620_CLKB;
 reg [1:16] _3I4365_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1310 (_3I4365_$1I4488_$1I4620_CLKB, _3I4365_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _3I4365_$1I4488_$1I4620_DIA;
 reg [1:16] _3I4365_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1311_7 (_3I4365_$1I4488_$1I4620_DIA[7], _3I4365_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1311_6 (_3I4365_$1I4488_$1I4620_DIA[6], _3I4365_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1311_5 (_3I4365_$1I4488_$1I4620_DIA[5], _3I4365_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1311_4 (_3I4365_$1I4488_$1I4620_DIA[4], _3I4365_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1311_3 (_3I4365_$1I4488_$1I4620_DIA[3], _3I4365_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1311_2 (_3I4365_$1I4488_$1I4620_DIA[2], _3I4365_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1311_1 (_3I4365_$1I4488_$1I4620_DIA[1], _3I4365_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1311_0 (_3I4365_$1I4488_$1I4620_DIA[0], _3I4365_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _3I4365_$1I4488_$1I4620_DIB;
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1312_15 (_3I4365_$1I4488_$1I4620_DIB[15], _3I4365_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1312_14 (_3I4365_$1I4488_$1I4620_DIB[14], _3I4365_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1312_13 (_3I4365_$1I4488_$1I4620_DIB[13], _3I4365_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1312_12 (_3I4365_$1I4488_$1I4620_DIB[12], _3I4365_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1312_11 (_3I4365_$1I4488_$1I4620_DIB[11], _3I4365_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1312_10 (_3I4365_$1I4488_$1I4620_DIB[10], _3I4365_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1312_9 (_3I4365_$1I4488_$1I4620_DIB[9], _3I4365_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1312_8 (_3I4365_$1I4488_$1I4620_DIB[8], _3I4365_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1312_7 (_3I4365_$1I4488_$1I4620_DIB[7], _3I4365_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1312_6 (_3I4365_$1I4488_$1I4620_DIB[6], _3I4365_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1312_5 (_3I4365_$1I4488_$1I4620_DIB[5], _3I4365_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1312_4 (_3I4365_$1I4488_$1I4620_DIB[4], _3I4365_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1312_3 (_3I4365_$1I4488_$1I4620_DIB[3], _3I4365_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1312_2 (_3I4365_$1I4488_$1I4620_DIB[2], _3I4365_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1312_1 (_3I4365_$1I4488_$1I4620_DIB[1], _3I4365_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1312_0 (_3I4365_$1I4488_$1I4620_DIB[0], _3I4365_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _3I4365_$1I4488_$1I4620_DIPA;
 reg [1:16] _3I4365_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1313_0 (_3I4365_$1I4488_$1I4620_DIPA[0], _3I4365_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _3I4365_$1I4488_$1I4620_DIPB;
 reg [1:16] _3I4365_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1314_1 (_3I4365_$1I4488_$1I4620_DIPB[1], _3I4365_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _3I4365_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1314_0 (_3I4365_$1I4488_$1I4620_DIPB[0], _3I4365_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _3I4365_$1I4488_$1I4620_ENA;
 reg [1:16] _3I4365_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1315 (_3I4365_$1I4488_$1I4620_ENA, _3I4365_$1I4488_$1I4620_ENA__vlIN);

 wire  _3I4365_$1I4488_$1I4620_ENB;
 reg [1:16] _3I4365_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1316 (_3I4365_$1I4488_$1I4620_ENB, _3I4365_$1I4488_$1I4620_ENB__vlIN);

 wire  _3I4365_$1I4488_$1I4620_SSRA;
 reg [1:16] _3I4365_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1317 (_3I4365_$1I4488_$1I4620_SSRA, _3I4365_$1I4488_$1I4620_SSRA__vlIN);

 wire  _3I4365_$1I4488_$1I4620_SSRB;
 reg [1:16] _3I4365_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1318 (_3I4365_$1I4488_$1I4620_SSRB, _3I4365_$1I4488_$1I4620_SSRB__vlIN);

 wire  _3I4365_$1I4488_$1I4620_WEA;
 reg [1:16] _3I4365_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1319 (_3I4365_$1I4488_$1I4620_WEA, _3I4365_$1I4488_$1I4620_WEA__vlIN);

 wire  _3I4365_$1I4488_$1I4620_WEB;
 reg [1:16] _3I4365_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1320 (_3I4365_$1I4488_$1I4620_WEB, _3I4365_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _3I4365_$1I4488_$1I4620 ( _3I4365_$1I4488_$1I4620_DOA , _3I4365_$1I4488_$1I4620_DOB , _3I4365_$1I4488_$1I4620_DOPA , _3I4365_$1I4488_$1I4620_DOPB , _3I4365_$1I4488_$1I4620_ADDRA , _3I4365_$1I4488_$1I4620_ADDRB , _3I4365_$1I4488_$1I4620_CLKA , _3I4365_$1I4488_$1I4620_CLKB , _3I4365_$1I4488_$1I4620_DIA , _3I4365_$1I4488_$1I4620_DIB , _3I4365_$1I4488_$1I4620_DIPA , _3I4365_$1I4488_$1I4620_DIPB , _3I4365_$1I4488_$1I4620_ENA , _3I4365_$1I4488_$1I4620_ENB , _3I4365_$1I4488_$1I4620_SSRA , _3I4365_$1I4488_$1I4620_SSRB , _3I4365_$1I4488_$1I4620_WEA , _3I4365_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4329_$1I4488_$1I4621_DOA;

 wire [15:0] _3I4329_$1I4488_$1I4621_DOB;

 wire [0:0] _3I4329_$1I4488_$1I4621_DOPA;

 wire [1:0] _3I4329_$1I4488_$1I4621_DOPB;

 wire [10:0] _3I4329_$1I4488_$1I4621_ADDRA;
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1321_10 (_3I4329_$1I4488_$1I4621_ADDRA[10], _3I4329_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1321_9 (_3I4329_$1I4488_$1I4621_ADDRA[9], _3I4329_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1321_8 (_3I4329_$1I4488_$1I4621_ADDRA[8], _3I4329_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1321_7 (_3I4329_$1I4488_$1I4621_ADDRA[7], _3I4329_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1321_6 (_3I4329_$1I4488_$1I4621_ADDRA[6], _3I4329_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1321_5 (_3I4329_$1I4488_$1I4621_ADDRA[5], _3I4329_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1321_4 (_3I4329_$1I4488_$1I4621_ADDRA[4], _3I4329_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1321_3 (_3I4329_$1I4488_$1I4621_ADDRA[3], _3I4329_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1321_2 (_3I4329_$1I4488_$1I4621_ADDRA[2], _3I4329_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1321_1 (_3I4329_$1I4488_$1I4621_ADDRA[1], _3I4329_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1321_0 (_3I4329_$1I4488_$1I4621_ADDRA[0], _3I4329_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _3I4329_$1I4488_$1I4621_ADDRB;
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_1322_9 (_3I4329_$1I4488_$1I4621_ADDRB[9], _3I4329_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_1322_8 (_3I4329_$1I4488_$1I4621_ADDRB[8], _3I4329_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_1322_7 (_3I4329_$1I4488_$1I4621_ADDRB[7], _3I4329_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_1322_6 (_3I4329_$1I4488_$1I4621_ADDRB[6], _3I4329_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_1322_5 (_3I4329_$1I4488_$1I4621_ADDRB[5], _3I4329_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_1322_4 (_3I4329_$1I4488_$1I4621_ADDRB[4], _3I4329_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_1322_3 (_3I4329_$1I4488_$1I4621_ADDRB[3], _3I4329_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_1322_2 (_3I4329_$1I4488_$1I4621_ADDRB[2], _3I4329_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_1322_1 (_3I4329_$1I4488_$1I4621_ADDRB[1], _3I4329_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_1322_0 (_3I4329_$1I4488_$1I4621_ADDRB[0], _3I4329_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _3I4329_$1I4488_$1I4621_CLKA;
 reg [1:16] _3I4329_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_1323 (_3I4329_$1I4488_$1I4621_CLKA, _3I4329_$1I4488_$1I4621_CLKA__vlIN);

 wire  _3I4329_$1I4488_$1I4621_CLKB;
 reg [1:16] _3I4329_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_1324 (_3I4329_$1I4488_$1I4621_CLKB, _3I4329_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _3I4329_$1I4488_$1I4621_DIA;
 reg [1:16] _3I4329_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_1325_7 (_3I4329_$1I4488_$1I4621_DIA[7], _3I4329_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_1325_6 (_3I4329_$1I4488_$1I4621_DIA[6], _3I4329_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_1325_5 (_3I4329_$1I4488_$1I4621_DIA[5], _3I4329_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_1325_4 (_3I4329_$1I4488_$1I4621_DIA[4], _3I4329_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_1325_3 (_3I4329_$1I4488_$1I4621_DIA[3], _3I4329_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_1325_2 (_3I4329_$1I4488_$1I4621_DIA[2], _3I4329_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_1325_1 (_3I4329_$1I4488_$1I4621_DIA[1], _3I4329_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_1325_0 (_3I4329_$1I4488_$1I4621_DIA[0], _3I4329_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _3I4329_$1I4488_$1I4621_DIB;
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_1326_15 (_3I4329_$1I4488_$1I4621_DIB[15], _3I4329_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_1326_14 (_3I4329_$1I4488_$1I4621_DIB[14], _3I4329_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_1326_13 (_3I4329_$1I4488_$1I4621_DIB[13], _3I4329_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_1326_12 (_3I4329_$1I4488_$1I4621_DIB[12], _3I4329_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_1326_11 (_3I4329_$1I4488_$1I4621_DIB[11], _3I4329_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_1326_10 (_3I4329_$1I4488_$1I4621_DIB[10], _3I4329_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_1326_9 (_3I4329_$1I4488_$1I4621_DIB[9], _3I4329_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_1326_8 (_3I4329_$1I4488_$1I4621_DIB[8], _3I4329_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_1326_7 (_3I4329_$1I4488_$1I4621_DIB[7], _3I4329_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_1326_6 (_3I4329_$1I4488_$1I4621_DIB[6], _3I4329_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_1326_5 (_3I4329_$1I4488_$1I4621_DIB[5], _3I4329_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_1326_4 (_3I4329_$1I4488_$1I4621_DIB[4], _3I4329_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_1326_3 (_3I4329_$1I4488_$1I4621_DIB[3], _3I4329_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_1326_2 (_3I4329_$1I4488_$1I4621_DIB[2], _3I4329_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_1326_1 (_3I4329_$1I4488_$1I4621_DIB[1], _3I4329_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_1326_0 (_3I4329_$1I4488_$1I4621_DIB[0], _3I4329_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _3I4329_$1I4488_$1I4621_DIPA;
 reg [1:16] _3I4329_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_1327_0 (_3I4329_$1I4488_$1I4621_DIPA[0], _3I4329_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _3I4329_$1I4488_$1I4621_DIPB;
 reg [1:16] _3I4329_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_1328_1 (_3I4329_$1I4488_$1I4621_DIPB[1], _3I4329_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_1328_0 (_3I4329_$1I4488_$1I4621_DIPB[0], _3I4329_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _3I4329_$1I4488_$1I4621_ENA;
 reg [1:16] _3I4329_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_1329 (_3I4329_$1I4488_$1I4621_ENA, _3I4329_$1I4488_$1I4621_ENA__vlIN);

 wire  _3I4329_$1I4488_$1I4621_ENB;
 reg [1:16] _3I4329_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_1330 (_3I4329_$1I4488_$1I4621_ENB, _3I4329_$1I4488_$1I4621_ENB__vlIN);

 wire  _3I4329_$1I4488_$1I4621_SSRA;
 reg [1:16] _3I4329_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_1331 (_3I4329_$1I4488_$1I4621_SSRA, _3I4329_$1I4488_$1I4621_SSRA__vlIN);

 wire  _3I4329_$1I4488_$1I4621_SSRB;
 reg [1:16] _3I4329_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_1332 (_3I4329_$1I4488_$1I4621_SSRB, _3I4329_$1I4488_$1I4621_SSRB__vlIN);

 wire  _3I4329_$1I4488_$1I4621_WEA;
 reg [1:16] _3I4329_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_1333 (_3I4329_$1I4488_$1I4621_WEA, _3I4329_$1I4488_$1I4621_WEA__vlIN);

 wire  _3I4329_$1I4488_$1I4621_WEB;
 reg [1:16] _3I4329_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_1334 (_3I4329_$1I4488_$1I4621_WEB, _3I4329_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _3I4329_$1I4488_$1I4621 ( _3I4329_$1I4488_$1I4621_DOA , _3I4329_$1I4488_$1I4621_DOB , _3I4329_$1I4488_$1I4621_DOPA , _3I4329_$1I4488_$1I4621_DOPB , _3I4329_$1I4488_$1I4621_ADDRA , _3I4329_$1I4488_$1I4621_ADDRB , _3I4329_$1I4488_$1I4621_CLKA , _3I4329_$1I4488_$1I4621_CLKB , _3I4329_$1I4488_$1I4621_DIA , _3I4329_$1I4488_$1I4621_DIB , _3I4329_$1I4488_$1I4621_DIPA , _3I4329_$1I4488_$1I4621_DIPB , _3I4329_$1I4488_$1I4621_ENA , _3I4329_$1I4488_$1I4621_ENB , _3I4329_$1I4488_$1I4621_SSRA , _3I4329_$1I4488_$1I4621_SSRB , _3I4329_$1I4488_$1I4621_WEA , _3I4329_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _3I4329_$1I4488_$1I4620_DOA;

 wire [15:0] _3I4329_$1I4488_$1I4620_DOB;

 wire [0:0] _3I4329_$1I4488_$1I4620_DOPA;

 wire [1:0] _3I4329_$1I4488_$1I4620_DOPB;

 wire [10:0] _3I4329_$1I4488_$1I4620_ADDRA;
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_1335_10 (_3I4329_$1I4488_$1I4620_ADDRA[10], _3I4329_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_1335_9 (_3I4329_$1I4488_$1I4620_ADDRA[9], _3I4329_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_1335_8 (_3I4329_$1I4488_$1I4620_ADDRA[8], _3I4329_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_1335_7 (_3I4329_$1I4488_$1I4620_ADDRA[7], _3I4329_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_1335_6 (_3I4329_$1I4488_$1I4620_ADDRA[6], _3I4329_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_1335_5 (_3I4329_$1I4488_$1I4620_ADDRA[5], _3I4329_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_1335_4 (_3I4329_$1I4488_$1I4620_ADDRA[4], _3I4329_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_1335_3 (_3I4329_$1I4488_$1I4620_ADDRA[3], _3I4329_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_1335_2 (_3I4329_$1I4488_$1I4620_ADDRA[2], _3I4329_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_1335_1 (_3I4329_$1I4488_$1I4620_ADDRA[1], _3I4329_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_1335_0 (_3I4329_$1I4488_$1I4620_ADDRA[0], _3I4329_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _3I4329_$1I4488_$1I4620_ADDRB;
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1336_9 (_3I4329_$1I4488_$1I4620_ADDRB[9], _3I4329_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1336_8 (_3I4329_$1I4488_$1I4620_ADDRB[8], _3I4329_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1336_7 (_3I4329_$1I4488_$1I4620_ADDRB[7], _3I4329_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1336_6 (_3I4329_$1I4488_$1I4620_ADDRB[6], _3I4329_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1336_5 (_3I4329_$1I4488_$1I4620_ADDRB[5], _3I4329_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1336_4 (_3I4329_$1I4488_$1I4620_ADDRB[4], _3I4329_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1336_3 (_3I4329_$1I4488_$1I4620_ADDRB[3], _3I4329_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1336_2 (_3I4329_$1I4488_$1I4620_ADDRB[2], _3I4329_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1336_1 (_3I4329_$1I4488_$1I4620_ADDRB[1], _3I4329_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1336_0 (_3I4329_$1I4488_$1I4620_ADDRB[0], _3I4329_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _3I4329_$1I4488_$1I4620_CLKA;
 reg [1:16] _3I4329_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1337 (_3I4329_$1I4488_$1I4620_CLKA, _3I4329_$1I4488_$1I4620_CLKA__vlIN);

 wire  _3I4329_$1I4488_$1I4620_CLKB;
 reg [1:16] _3I4329_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1338 (_3I4329_$1I4488_$1I4620_CLKB, _3I4329_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _3I4329_$1I4488_$1I4620_DIA;
 reg [1:16] _3I4329_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1339_7 (_3I4329_$1I4488_$1I4620_DIA[7], _3I4329_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1339_6 (_3I4329_$1I4488_$1I4620_DIA[6], _3I4329_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1339_5 (_3I4329_$1I4488_$1I4620_DIA[5], _3I4329_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1339_4 (_3I4329_$1I4488_$1I4620_DIA[4], _3I4329_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1339_3 (_3I4329_$1I4488_$1I4620_DIA[3], _3I4329_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1339_2 (_3I4329_$1I4488_$1I4620_DIA[2], _3I4329_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1339_1 (_3I4329_$1I4488_$1I4620_DIA[1], _3I4329_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1339_0 (_3I4329_$1I4488_$1I4620_DIA[0], _3I4329_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _3I4329_$1I4488_$1I4620_DIB;
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1340_15 (_3I4329_$1I4488_$1I4620_DIB[15], _3I4329_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1340_14 (_3I4329_$1I4488_$1I4620_DIB[14], _3I4329_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1340_13 (_3I4329_$1I4488_$1I4620_DIB[13], _3I4329_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1340_12 (_3I4329_$1I4488_$1I4620_DIB[12], _3I4329_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1340_11 (_3I4329_$1I4488_$1I4620_DIB[11], _3I4329_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1340_10 (_3I4329_$1I4488_$1I4620_DIB[10], _3I4329_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1340_9 (_3I4329_$1I4488_$1I4620_DIB[9], _3I4329_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1340_8 (_3I4329_$1I4488_$1I4620_DIB[8], _3I4329_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1340_7 (_3I4329_$1I4488_$1I4620_DIB[7], _3I4329_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1340_6 (_3I4329_$1I4488_$1I4620_DIB[6], _3I4329_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1340_5 (_3I4329_$1I4488_$1I4620_DIB[5], _3I4329_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1340_4 (_3I4329_$1I4488_$1I4620_DIB[4], _3I4329_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1340_3 (_3I4329_$1I4488_$1I4620_DIB[3], _3I4329_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1340_2 (_3I4329_$1I4488_$1I4620_DIB[2], _3I4329_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1340_1 (_3I4329_$1I4488_$1I4620_DIB[1], _3I4329_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1340_0 (_3I4329_$1I4488_$1I4620_DIB[0], _3I4329_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _3I4329_$1I4488_$1I4620_DIPA;
 reg [1:16] _3I4329_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1341_0 (_3I4329_$1I4488_$1I4620_DIPA[0], _3I4329_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _3I4329_$1I4488_$1I4620_DIPB;
 reg [1:16] _3I4329_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1342_1 (_3I4329_$1I4488_$1I4620_DIPB[1], _3I4329_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _3I4329_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1342_0 (_3I4329_$1I4488_$1I4620_DIPB[0], _3I4329_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _3I4329_$1I4488_$1I4620_ENA;
 reg [1:16] _3I4329_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1343 (_3I4329_$1I4488_$1I4620_ENA, _3I4329_$1I4488_$1I4620_ENA__vlIN);

 wire  _3I4329_$1I4488_$1I4620_ENB;
 reg [1:16] _3I4329_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1344 (_3I4329_$1I4488_$1I4620_ENB, _3I4329_$1I4488_$1I4620_ENB__vlIN);

 wire  _3I4329_$1I4488_$1I4620_SSRA;
 reg [1:16] _3I4329_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1345 (_3I4329_$1I4488_$1I4620_SSRA, _3I4329_$1I4488_$1I4620_SSRA__vlIN);

 wire  _3I4329_$1I4488_$1I4620_SSRB;
 reg [1:16] _3I4329_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1346 (_3I4329_$1I4488_$1I4620_SSRB, _3I4329_$1I4488_$1I4620_SSRB__vlIN);

 wire  _3I4329_$1I4488_$1I4620_WEA;
 reg [1:16] _3I4329_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1347 (_3I4329_$1I4488_$1I4620_WEA, _3I4329_$1I4488_$1I4620_WEA__vlIN);

 wire  _3I4329_$1I4488_$1I4620_WEB;
 reg [1:16] _3I4329_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1348 (_3I4329_$1I4488_$1I4620_WEB, _3I4329_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _3I4329_$1I4488_$1I4620 ( _3I4329_$1I4488_$1I4620_DOA , _3I4329_$1I4488_$1I4620_DOB , _3I4329_$1I4488_$1I4620_DOPA , _3I4329_$1I4488_$1I4620_DOPB , _3I4329_$1I4488_$1I4620_ADDRA , _3I4329_$1I4488_$1I4620_ADDRB , _3I4329_$1I4488_$1I4620_CLKA , _3I4329_$1I4488_$1I4620_CLKB , _3I4329_$1I4488_$1I4620_DIA , _3I4329_$1I4488_$1I4620_DIB , _3I4329_$1I4488_$1I4620_DIPA , _3I4329_$1I4488_$1I4620_DIPB , _3I4329_$1I4488_$1I4620_ENA , _3I4329_$1I4488_$1I4620_ENB , _3I4329_$1I4488_$1I4620_SSRA , _3I4329_$1I4488_$1I4620_SSRB , _3I4329_$1I4488_$1I4620_WEA , _3I4329_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [4:0] _3I4274_$1I4152_din;
 reg [1:16] _3I4274_$1I4152_din_4__vlIN;
 cstw cstw_1349_4 (_3I4274_$1I4152_din[4], _3I4274_$1I4152_din_4__vlIN);
 reg [1:16] _3I4274_$1I4152_din_3__vlIN;
 cstw cstw_1349_3 (_3I4274_$1I4152_din[3], _3I4274_$1I4152_din_3__vlIN);
 reg [1:16] _3I4274_$1I4152_din_2__vlIN;
 cstw cstw_1349_2 (_3I4274_$1I4152_din[2], _3I4274_$1I4152_din_2__vlIN);
 reg [1:16] _3I4274_$1I4152_din_1__vlIN;
 cstw cstw_1349_1 (_3I4274_$1I4152_din[1], _3I4274_$1I4152_din_1__vlIN);
 reg [1:16] _3I4274_$1I4152_din_0__vlIN;
 cstw cstw_1349_0 (_3I4274_$1I4152_din[0], _3I4274_$1I4152_din_0__vlIN);

 wire  _3I4274_$1I4152_wr_en;
 reg [1:16] _3I4274_$1I4152_wr_en__vlIN;
 cstw cstw_1350 (_3I4274_$1I4152_wr_en, _3I4274_$1I4152_wr_en__vlIN);

 wire  _3I4274_$1I4152_wr_clk;
 reg [1:16] _3I4274_$1I4152_wr_clk__vlIN;
 cstw cstw_1351 (_3I4274_$1I4152_wr_clk, _3I4274_$1I4152_wr_clk__vlIN);

 wire  _3I4274_$1I4152_rd_en;
 reg [1:16] _3I4274_$1I4152_rd_en__vlIN;
 cstw cstw_1352 (_3I4274_$1I4152_rd_en, _3I4274_$1I4152_rd_en__vlIN);

 wire  _3I4274_$1I4152_rd_clk;
 reg [1:16] _3I4274_$1I4152_rd_clk__vlIN;
 cstw cstw_1353 (_3I4274_$1I4152_rd_clk, _3I4274_$1I4152_rd_clk__vlIN);

 wire  _3I4274_$1I4152_ainit;
 reg [1:16] _3I4274_$1I4152_ainit__vlIN;
 cstw cstw_1354 (_3I4274_$1I4152_ainit, _3I4274_$1I4152_ainit__vlIN);

 wire [4:0] _3I4274_$1I4152_dout;

 wire  _3I4274_$1I4152_full;

 wire  _3I4274_$1I4152_empty;

 af_clb_5x31rpm _3I4274_$1I4152 ( _3I4274_$1I4152_din , _3I4274_$1I4152_wr_en , _3I4274_$1I4152_wr_clk , _3I4274_$1I4152_rd_en , _3I4274_$1I4152_rd_clk , _3I4274_$1I4152_ainit , _3I4274_$1I4152_dout , _3I4274_$1I4152_full , _3I4274_$1I4152_empty  );

// ----------------------------------- //

 wire  _3I4274_$1I3863_CHBONDDONE;

 wire [3:0] _3I4274_$1I3863_CHBONDO;

 wire  _3I4274_$1I3863_CONFIGOUT;

 wire [1:0] _3I4274_$1I3863_RXBUFSTATUS;

 wire [3:0] _3I4274_$1I3863_RXCHARISCOMMA;

 wire [3:0] _3I4274_$1I3863_RXCHARISK;

 wire  _3I4274_$1I3863_RXCHECKINGCRC;

 wire [2:0] _3I4274_$1I3863_RXCLKCORCNT;

 wire  _3I4274_$1I3863_RXCOMMADET;

 wire  _3I4274_$1I3863_RXCRCERR;

 wire [31:0] _3I4274_$1I3863_RXDATA;

 wire [3:0] _3I4274_$1I3863_RXDISPERR;

 wire [1:0] _3I4274_$1I3863_RXLOSSOFSYNC;

 wire [3:0] _3I4274_$1I3863_RXNOTINTABLE;

 wire  _3I4274_$1I3863_RXREALIGN;

 wire  _3I4274_$1I3863_RXRECCLK;

 wire [3:0] _3I4274_$1I3863_RXRUNDISP;

 wire  _3I4274_$1I3863_TXBUFERR;

 wire [3:0] _3I4274_$1I3863_TXKERR;

 wire  _3I4274_$1I3863_TXN;

 wire  _3I4274_$1I3863_TXP;

 wire [3:0] _3I4274_$1I3863_TXRUNDISP;

 wire  _3I4274_$1I3863_BREFCLK;
 reg [1:16] _3I4274_$1I3863_BREFCLK__vlIN;
 cstw cstw_1355 (_3I4274_$1I3863_BREFCLK, _3I4274_$1I3863_BREFCLK__vlIN);

 wire  _3I4274_$1I3863_BREFCLK2;
 reg [1:16] _3I4274_$1I3863_BREFCLK2__vlIN;
 cstw cstw_1356 (_3I4274_$1I3863_BREFCLK2, _3I4274_$1I3863_BREFCLK2__vlIN);

 wire [3:0] _3I4274_$1I3863_CHBONDI;
 reg [1:16] _3I4274_$1I3863_CHBONDI_3__vlIN;
 cstw cstw_1357_3 (_3I4274_$1I3863_CHBONDI[3], _3I4274_$1I3863_CHBONDI_3__vlIN);
 reg [1:16] _3I4274_$1I3863_CHBONDI_2__vlIN;
 cstw cstw_1357_2 (_3I4274_$1I3863_CHBONDI[2], _3I4274_$1I3863_CHBONDI_2__vlIN);
 reg [1:16] _3I4274_$1I3863_CHBONDI_1__vlIN;
 cstw cstw_1357_1 (_3I4274_$1I3863_CHBONDI[1], _3I4274_$1I3863_CHBONDI_1__vlIN);
 reg [1:16] _3I4274_$1I3863_CHBONDI_0__vlIN;
 cstw cstw_1357_0 (_3I4274_$1I3863_CHBONDI[0], _3I4274_$1I3863_CHBONDI_0__vlIN);

 wire  _3I4274_$1I3863_CONFIGENABLE;
 reg [1:16] _3I4274_$1I3863_CONFIGENABLE__vlIN;
 cstw cstw_1358 (_3I4274_$1I3863_CONFIGENABLE, _3I4274_$1I3863_CONFIGENABLE__vlIN);

 wire  _3I4274_$1I3863_CONFIGIN;
 reg [1:16] _3I4274_$1I3863_CONFIGIN__vlIN;
 cstw cstw_1359 (_3I4274_$1I3863_CONFIGIN, _3I4274_$1I3863_CONFIGIN__vlIN);

 wire  _3I4274_$1I3863_ENCHANSYNC;
 reg [1:16] _3I4274_$1I3863_ENCHANSYNC__vlIN;
 cstw cstw_1360 (_3I4274_$1I3863_ENCHANSYNC, _3I4274_$1I3863_ENCHANSYNC__vlIN);

 wire  _3I4274_$1I3863_ENMCOMMAALIGN;
 reg [1:16] _3I4274_$1I3863_ENMCOMMAALIGN__vlIN;
 cstw cstw_1361 (_3I4274_$1I3863_ENMCOMMAALIGN, _3I4274_$1I3863_ENMCOMMAALIGN__vlIN);

 wire  _3I4274_$1I3863_ENPCOMMAALIGN;
 reg [1:16] _3I4274_$1I3863_ENPCOMMAALIGN__vlIN;
 cstw cstw_1362 (_3I4274_$1I3863_ENPCOMMAALIGN, _3I4274_$1I3863_ENPCOMMAALIGN__vlIN);

 wire [1:0] _3I4274_$1I3863_LOOPBACK;
 reg [1:16] _3I4274_$1I3863_LOOPBACK_1__vlIN;
 cstw cstw_1363_1 (_3I4274_$1I3863_LOOPBACK[1], _3I4274_$1I3863_LOOPBACK_1__vlIN);
 reg [1:16] _3I4274_$1I3863_LOOPBACK_0__vlIN;
 cstw cstw_1363_0 (_3I4274_$1I3863_LOOPBACK[0], _3I4274_$1I3863_LOOPBACK_0__vlIN);

 wire  _3I4274_$1I3863_POWERDOWN;
 reg [1:16] _3I4274_$1I3863_POWERDOWN__vlIN;
 cstw cstw_1364 (_3I4274_$1I3863_POWERDOWN, _3I4274_$1I3863_POWERDOWN__vlIN);

 wire  _3I4274_$1I3863_REFCLK;
 reg [1:16] _3I4274_$1I3863_REFCLK__vlIN;
 cstw cstw_1365 (_3I4274_$1I3863_REFCLK, _3I4274_$1I3863_REFCLK__vlIN);

 wire  _3I4274_$1I3863_REFCLK2;
 reg [1:16] _3I4274_$1I3863_REFCLK2__vlIN;
 cstw cstw_1366 (_3I4274_$1I3863_REFCLK2, _3I4274_$1I3863_REFCLK2__vlIN);

 wire  _3I4274_$1I3863_REFCLKSEL;
 reg [1:16] _3I4274_$1I3863_REFCLKSEL__vlIN;
 cstw cstw_1367 (_3I4274_$1I3863_REFCLKSEL, _3I4274_$1I3863_REFCLKSEL__vlIN);

 wire  _3I4274_$1I3863_RXN;
 reg [1:16] _3I4274_$1I3863_RXN__vlIN;
 cstw cstw_1368 (_3I4274_$1I3863_RXN, _3I4274_$1I3863_RXN__vlIN);

 wire  _3I4274_$1I3863_RXP;
 reg [1:16] _3I4274_$1I3863_RXP__vlIN;
 cstw cstw_1369 (_3I4274_$1I3863_RXP, _3I4274_$1I3863_RXP__vlIN);

 wire  _3I4274_$1I3863_RXPOLARITY;
 reg [1:16] _3I4274_$1I3863_RXPOLARITY__vlIN;
 cstw cstw_1370 (_3I4274_$1I3863_RXPOLARITY, _3I4274_$1I3863_RXPOLARITY__vlIN);

 wire  _3I4274_$1I3863_RXRESET;
 reg [1:16] _3I4274_$1I3863_RXRESET__vlIN;
 cstw cstw_1371 (_3I4274_$1I3863_RXRESET, _3I4274_$1I3863_RXRESET__vlIN);

 wire  _3I4274_$1I3863_RXUSRCLK;
 reg [1:16] _3I4274_$1I3863_RXUSRCLK__vlIN;
 cstw cstw_1372 (_3I4274_$1I3863_RXUSRCLK, _3I4274_$1I3863_RXUSRCLK__vlIN);

 wire  _3I4274_$1I3863_RXUSRCLK2;
 reg [1:16] _3I4274_$1I3863_RXUSRCLK2__vlIN;
 cstw cstw_1373 (_3I4274_$1I3863_RXUSRCLK2, _3I4274_$1I3863_RXUSRCLK2__vlIN);

 wire [3:0] _3I4274_$1I3863_TXBYPASS8B10B;
 reg [1:16] _3I4274_$1I3863_TXBYPASS8B10B_3__vlIN;
 cstw cstw_1374_3 (_3I4274_$1I3863_TXBYPASS8B10B[3], _3I4274_$1I3863_TXBYPASS8B10B_3__vlIN);
 reg [1:16] _3I4274_$1I3863_TXBYPASS8B10B_2__vlIN;
 cstw cstw_1374_2 (_3I4274_$1I3863_TXBYPASS8B10B[2], _3I4274_$1I3863_TXBYPASS8B10B_2__vlIN);
 reg [1:16] _3I4274_$1I3863_TXBYPASS8B10B_1__vlIN;
 cstw cstw_1374_1 (_3I4274_$1I3863_TXBYPASS8B10B[1], _3I4274_$1I3863_TXBYPASS8B10B_1__vlIN);
 reg [1:16] _3I4274_$1I3863_TXBYPASS8B10B_0__vlIN;
 cstw cstw_1374_0 (_3I4274_$1I3863_TXBYPASS8B10B[0], _3I4274_$1I3863_TXBYPASS8B10B_0__vlIN);

 wire [3:0] _3I4274_$1I3863_TXCHARDISPMODE;
 reg [1:16] _3I4274_$1I3863_TXCHARDISPMODE_3__vlIN;
 cstw cstw_1375_3 (_3I4274_$1I3863_TXCHARDISPMODE[3], _3I4274_$1I3863_TXCHARDISPMODE_3__vlIN);
 reg [1:16] _3I4274_$1I3863_TXCHARDISPMODE_2__vlIN;
 cstw cstw_1375_2 (_3I4274_$1I3863_TXCHARDISPMODE[2], _3I4274_$1I3863_TXCHARDISPMODE_2__vlIN);
 reg [1:16] _3I4274_$1I3863_TXCHARDISPMODE_1__vlIN;
 cstw cstw_1375_1 (_3I4274_$1I3863_TXCHARDISPMODE[1], _3I4274_$1I3863_TXCHARDISPMODE_1__vlIN);
 reg [1:16] _3I4274_$1I3863_TXCHARDISPMODE_0__vlIN;
 cstw cstw_1375_0 (_3I4274_$1I3863_TXCHARDISPMODE[0], _3I4274_$1I3863_TXCHARDISPMODE_0__vlIN);

 wire [3:0] _3I4274_$1I3863_TXCHARDISPVAL;
 reg [1:16] _3I4274_$1I3863_TXCHARDISPVAL_3__vlIN;
 cstw cstw_1376_3 (_3I4274_$1I3863_TXCHARDISPVAL[3], _3I4274_$1I3863_TXCHARDISPVAL_3__vlIN);
 reg [1:16] _3I4274_$1I3863_TXCHARDISPVAL_2__vlIN;
 cstw cstw_1376_2 (_3I4274_$1I3863_TXCHARDISPVAL[2], _3I4274_$1I3863_TXCHARDISPVAL_2__vlIN);
 reg [1:16] _3I4274_$1I3863_TXCHARDISPVAL_1__vlIN;
 cstw cstw_1376_1 (_3I4274_$1I3863_TXCHARDISPVAL[1], _3I4274_$1I3863_TXCHARDISPVAL_1__vlIN);
 reg [1:16] _3I4274_$1I3863_TXCHARDISPVAL_0__vlIN;
 cstw cstw_1376_0 (_3I4274_$1I3863_TXCHARDISPVAL[0], _3I4274_$1I3863_TXCHARDISPVAL_0__vlIN);

 wire [3:0] _3I4274_$1I3863_TXCHARISK;
 reg [1:16] _3I4274_$1I3863_TXCHARISK_3__vlIN;
 cstw cstw_1377_3 (_3I4274_$1I3863_TXCHARISK[3], _3I4274_$1I3863_TXCHARISK_3__vlIN);
 reg [1:16] _3I4274_$1I3863_TXCHARISK_2__vlIN;
 cstw cstw_1377_2 (_3I4274_$1I3863_TXCHARISK[2], _3I4274_$1I3863_TXCHARISK_2__vlIN);
 reg [1:16] _3I4274_$1I3863_TXCHARISK_1__vlIN;
 cstw cstw_1377_1 (_3I4274_$1I3863_TXCHARISK[1], _3I4274_$1I3863_TXCHARISK_1__vlIN);
 reg [1:16] _3I4274_$1I3863_TXCHARISK_0__vlIN;
 cstw cstw_1377_0 (_3I4274_$1I3863_TXCHARISK[0], _3I4274_$1I3863_TXCHARISK_0__vlIN);

 wire [31:0] _3I4274_$1I3863_TXDATA;
 reg [1:16] _3I4274_$1I3863_TXDATA_31__vlIN;
 cstw cstw_1378_31 (_3I4274_$1I3863_TXDATA[31], _3I4274_$1I3863_TXDATA_31__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_30__vlIN;
 cstw cstw_1378_30 (_3I4274_$1I3863_TXDATA[30], _3I4274_$1I3863_TXDATA_30__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_29__vlIN;
 cstw cstw_1378_29 (_3I4274_$1I3863_TXDATA[29], _3I4274_$1I3863_TXDATA_29__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_28__vlIN;
 cstw cstw_1378_28 (_3I4274_$1I3863_TXDATA[28], _3I4274_$1I3863_TXDATA_28__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_27__vlIN;
 cstw cstw_1378_27 (_3I4274_$1I3863_TXDATA[27], _3I4274_$1I3863_TXDATA_27__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_26__vlIN;
 cstw cstw_1378_26 (_3I4274_$1I3863_TXDATA[26], _3I4274_$1I3863_TXDATA_26__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_25__vlIN;
 cstw cstw_1378_25 (_3I4274_$1I3863_TXDATA[25], _3I4274_$1I3863_TXDATA_25__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_24__vlIN;
 cstw cstw_1378_24 (_3I4274_$1I3863_TXDATA[24], _3I4274_$1I3863_TXDATA_24__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_23__vlIN;
 cstw cstw_1378_23 (_3I4274_$1I3863_TXDATA[23], _3I4274_$1I3863_TXDATA_23__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_22__vlIN;
 cstw cstw_1378_22 (_3I4274_$1I3863_TXDATA[22], _3I4274_$1I3863_TXDATA_22__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_21__vlIN;
 cstw cstw_1378_21 (_3I4274_$1I3863_TXDATA[21], _3I4274_$1I3863_TXDATA_21__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_20__vlIN;
 cstw cstw_1378_20 (_3I4274_$1I3863_TXDATA[20], _3I4274_$1I3863_TXDATA_20__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_19__vlIN;
 cstw cstw_1378_19 (_3I4274_$1I3863_TXDATA[19], _3I4274_$1I3863_TXDATA_19__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_18__vlIN;
 cstw cstw_1378_18 (_3I4274_$1I3863_TXDATA[18], _3I4274_$1I3863_TXDATA_18__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_17__vlIN;
 cstw cstw_1378_17 (_3I4274_$1I3863_TXDATA[17], _3I4274_$1I3863_TXDATA_17__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_16__vlIN;
 cstw cstw_1378_16 (_3I4274_$1I3863_TXDATA[16], _3I4274_$1I3863_TXDATA_16__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_15__vlIN;
 cstw cstw_1378_15 (_3I4274_$1I3863_TXDATA[15], _3I4274_$1I3863_TXDATA_15__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_14__vlIN;
 cstw cstw_1378_14 (_3I4274_$1I3863_TXDATA[14], _3I4274_$1I3863_TXDATA_14__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_13__vlIN;
 cstw cstw_1378_13 (_3I4274_$1I3863_TXDATA[13], _3I4274_$1I3863_TXDATA_13__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_12__vlIN;
 cstw cstw_1378_12 (_3I4274_$1I3863_TXDATA[12], _3I4274_$1I3863_TXDATA_12__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_11__vlIN;
 cstw cstw_1378_11 (_3I4274_$1I3863_TXDATA[11], _3I4274_$1I3863_TXDATA_11__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_10__vlIN;
 cstw cstw_1378_10 (_3I4274_$1I3863_TXDATA[10], _3I4274_$1I3863_TXDATA_10__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_9__vlIN;
 cstw cstw_1378_9 (_3I4274_$1I3863_TXDATA[9], _3I4274_$1I3863_TXDATA_9__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_8__vlIN;
 cstw cstw_1378_8 (_3I4274_$1I3863_TXDATA[8], _3I4274_$1I3863_TXDATA_8__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_7__vlIN;
 cstw cstw_1378_7 (_3I4274_$1I3863_TXDATA[7], _3I4274_$1I3863_TXDATA_7__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_6__vlIN;
 cstw cstw_1378_6 (_3I4274_$1I3863_TXDATA[6], _3I4274_$1I3863_TXDATA_6__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_5__vlIN;
 cstw cstw_1378_5 (_3I4274_$1I3863_TXDATA[5], _3I4274_$1I3863_TXDATA_5__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_4__vlIN;
 cstw cstw_1378_4 (_3I4274_$1I3863_TXDATA[4], _3I4274_$1I3863_TXDATA_4__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_3__vlIN;
 cstw cstw_1378_3 (_3I4274_$1I3863_TXDATA[3], _3I4274_$1I3863_TXDATA_3__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_2__vlIN;
 cstw cstw_1378_2 (_3I4274_$1I3863_TXDATA[2], _3I4274_$1I3863_TXDATA_2__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_1__vlIN;
 cstw cstw_1378_1 (_3I4274_$1I3863_TXDATA[1], _3I4274_$1I3863_TXDATA_1__vlIN);
 reg [1:16] _3I4274_$1I3863_TXDATA_0__vlIN;
 cstw cstw_1378_0 (_3I4274_$1I3863_TXDATA[0], _3I4274_$1I3863_TXDATA_0__vlIN);

 wire  _3I4274_$1I3863_TXFORCECRCERR;
 reg [1:16] _3I4274_$1I3863_TXFORCECRCERR__vlIN;
 cstw cstw_1379 (_3I4274_$1I3863_TXFORCECRCERR, _3I4274_$1I3863_TXFORCECRCERR__vlIN);

 wire  _3I4274_$1I3863_TXINHIBIT;
 reg [1:16] _3I4274_$1I3863_TXINHIBIT__vlIN;
 cstw cstw_1380 (_3I4274_$1I3863_TXINHIBIT, _3I4274_$1I3863_TXINHIBIT__vlIN);

 wire  _3I4274_$1I3863_TXPOLARITY;
 reg [1:16] _3I4274_$1I3863_TXPOLARITY__vlIN;
 cstw cstw_1381 (_3I4274_$1I3863_TXPOLARITY, _3I4274_$1I3863_TXPOLARITY__vlIN);

 wire  _3I4274_$1I3863_TXRESET;
 reg [1:16] _3I4274_$1I3863_TXRESET__vlIN;
 cstw cstw_1382 (_3I4274_$1I3863_TXRESET, _3I4274_$1I3863_TXRESET__vlIN);

 wire  _3I4274_$1I3863_TXUSRCLK;
 reg [1:16] _3I4274_$1I3863_TXUSRCLK__vlIN;
 cstw cstw_1383 (_3I4274_$1I3863_TXUSRCLK, _3I4274_$1I3863_TXUSRCLK__vlIN);

 wire  _3I4274_$1I3863_TXUSRCLK2;
 reg [1:16] _3I4274_$1I3863_TXUSRCLK2__vlIN;
 cstw cstw_1384 (_3I4274_$1I3863_TXUSRCLK2, _3I4274_$1I3863_TXUSRCLK2__vlIN);

 GT_CUSTOM _3I4274_$1I3863 ( _3I4274_$1I3863_CHBONDDONE , _3I4274_$1I3863_CHBONDO , _3I4274_$1I3863_CONFIGOUT , _3I4274_$1I3863_RXBUFSTATUS , _3I4274_$1I3863_RXCHARISCOMMA , _3I4274_$1I3863_RXCHARISK , _3I4274_$1I3863_RXCHECKINGCRC , _3I4274_$1I3863_RXCLKCORCNT , _3I4274_$1I3863_RXCOMMADET , _3I4274_$1I3863_RXCRCERR , _3I4274_$1I3863_RXDATA , _3I4274_$1I3863_RXDISPERR , _3I4274_$1I3863_RXLOSSOFSYNC , _3I4274_$1I3863_RXNOTINTABLE , _3I4274_$1I3863_RXREALIGN , _3I4274_$1I3863_RXRECCLK , _3I4274_$1I3863_RXRUNDISP , _3I4274_$1I3863_TXBUFERR , _3I4274_$1I3863_TXKERR , _3I4274_$1I3863_TXN , _3I4274_$1I3863_TXP , _3I4274_$1I3863_TXRUNDISP , _3I4274_$1I3863_BREFCLK , _3I4274_$1I3863_BREFCLK2 , _3I4274_$1I3863_CHBONDI , _3I4274_$1I3863_CONFIGENABLE , _3I4274_$1I3863_CONFIGIN , _3I4274_$1I3863_ENCHANSYNC , _3I4274_$1I3863_ENMCOMMAALIGN , _3I4274_$1I3863_ENPCOMMAALIGN , _3I4274_$1I3863_LOOPBACK , _3I4274_$1I3863_POWERDOWN , _3I4274_$1I3863_REFCLK , _3I4274_$1I3863_REFCLK2 , _3I4274_$1I3863_REFCLKSEL , _3I4274_$1I3863_RXN , _3I4274_$1I3863_RXP , _3I4274_$1I3863_RXPOLARITY , _3I4274_$1I3863_RXRESET , _3I4274_$1I3863_RXUSRCLK , _3I4274_$1I3863_RXUSRCLK2 , _3I4274_$1I3863_TXBYPASS8B10B , _3I4274_$1I3863_TXCHARDISPMODE , _3I4274_$1I3863_TXCHARDISPVAL , _3I4274_$1I3863_TXCHARISK , _3I4274_$1I3863_TXDATA , _3I4274_$1I3863_TXFORCECRCERR , _3I4274_$1I3863_TXINHIBIT , _3I4274_$1I3863_TXPOLARITY , _3I4274_$1I3863_TXRESET , _3I4274_$1I3863_TXUSRCLK , _3I4274_$1I3863_TXUSRCLK2  );

// ----------------------------------- //

 wire [4:0] _3I4243_$1I4152_din;
 reg [1:16] _3I4243_$1I4152_din_4__vlIN;
 cstw cstw_1385_4 (_3I4243_$1I4152_din[4], _3I4243_$1I4152_din_4__vlIN);
 reg [1:16] _3I4243_$1I4152_din_3__vlIN;
 cstw cstw_1385_3 (_3I4243_$1I4152_din[3], _3I4243_$1I4152_din_3__vlIN);
 reg [1:16] _3I4243_$1I4152_din_2__vlIN;
 cstw cstw_1385_2 (_3I4243_$1I4152_din[2], _3I4243_$1I4152_din_2__vlIN);
 reg [1:16] _3I4243_$1I4152_din_1__vlIN;
 cstw cstw_1385_1 (_3I4243_$1I4152_din[1], _3I4243_$1I4152_din_1__vlIN);
 reg [1:16] _3I4243_$1I4152_din_0__vlIN;
 cstw cstw_1385_0 (_3I4243_$1I4152_din[0], _3I4243_$1I4152_din_0__vlIN);

 wire  _3I4243_$1I4152_wr_en;
 reg [1:16] _3I4243_$1I4152_wr_en__vlIN;
 cstw cstw_1386 (_3I4243_$1I4152_wr_en, _3I4243_$1I4152_wr_en__vlIN);

 wire  _3I4243_$1I4152_wr_clk;
 reg [1:16] _3I4243_$1I4152_wr_clk__vlIN;
 cstw cstw_1387 (_3I4243_$1I4152_wr_clk, _3I4243_$1I4152_wr_clk__vlIN);

 wire  _3I4243_$1I4152_rd_en;
 reg [1:16] _3I4243_$1I4152_rd_en__vlIN;
 cstw cstw_1388 (_3I4243_$1I4152_rd_en, _3I4243_$1I4152_rd_en__vlIN);

 wire  _3I4243_$1I4152_rd_clk;
 reg [1:16] _3I4243_$1I4152_rd_clk__vlIN;
 cstw cstw_1389 (_3I4243_$1I4152_rd_clk, _3I4243_$1I4152_rd_clk__vlIN);

 wire  _3I4243_$1I4152_ainit;
 reg [1:16] _3I4243_$1I4152_ainit__vlIN;
 cstw cstw_1390 (_3I4243_$1I4152_ainit, _3I4243_$1I4152_ainit__vlIN);

 wire [4:0] _3I4243_$1I4152_dout;

 wire  _3I4243_$1I4152_full;

 wire  _3I4243_$1I4152_empty;

 af_clb_5x31rpm _3I4243_$1I4152 ( _3I4243_$1I4152_din , _3I4243_$1I4152_wr_en , _3I4243_$1I4152_wr_clk , _3I4243_$1I4152_rd_en , _3I4243_$1I4152_rd_clk , _3I4243_$1I4152_ainit , _3I4243_$1I4152_dout , _3I4243_$1I4152_full , _3I4243_$1I4152_empty  );

// ----------------------------------- //

 wire  _3I4243_$1I3863_CHBONDDONE;

 wire [3:0] _3I4243_$1I3863_CHBONDO;

 wire  _3I4243_$1I3863_CONFIGOUT;

 wire [1:0] _3I4243_$1I3863_RXBUFSTATUS;

 wire [3:0] _3I4243_$1I3863_RXCHARISCOMMA;

 wire [3:0] _3I4243_$1I3863_RXCHARISK;

 wire  _3I4243_$1I3863_RXCHECKINGCRC;

 wire [2:0] _3I4243_$1I3863_RXCLKCORCNT;

 wire  _3I4243_$1I3863_RXCOMMADET;

 wire  _3I4243_$1I3863_RXCRCERR;

 wire [31:0] _3I4243_$1I3863_RXDATA;

 wire [3:0] _3I4243_$1I3863_RXDISPERR;

 wire [1:0] _3I4243_$1I3863_RXLOSSOFSYNC;

 wire [3:0] _3I4243_$1I3863_RXNOTINTABLE;

 wire  _3I4243_$1I3863_RXREALIGN;

 wire  _3I4243_$1I3863_RXRECCLK;

 wire [3:0] _3I4243_$1I3863_RXRUNDISP;

 wire  _3I4243_$1I3863_TXBUFERR;

 wire [3:0] _3I4243_$1I3863_TXKERR;

 wire  _3I4243_$1I3863_TXN;

 wire  _3I4243_$1I3863_TXP;

 wire [3:0] _3I4243_$1I3863_TXRUNDISP;

 wire  _3I4243_$1I3863_BREFCLK;
 reg [1:16] _3I4243_$1I3863_BREFCLK__vlIN;
 cstw cstw_1391 (_3I4243_$1I3863_BREFCLK, _3I4243_$1I3863_BREFCLK__vlIN);

 wire  _3I4243_$1I3863_BREFCLK2;
 reg [1:16] _3I4243_$1I3863_BREFCLK2__vlIN;
 cstw cstw_1392 (_3I4243_$1I3863_BREFCLK2, _3I4243_$1I3863_BREFCLK2__vlIN);

 wire [3:0] _3I4243_$1I3863_CHBONDI;
 reg [1:16] _3I4243_$1I3863_CHBONDI_3__vlIN;
 cstw cstw_1393_3 (_3I4243_$1I3863_CHBONDI[3], _3I4243_$1I3863_CHBONDI_3__vlIN);
 reg [1:16] _3I4243_$1I3863_CHBONDI_2__vlIN;
 cstw cstw_1393_2 (_3I4243_$1I3863_CHBONDI[2], _3I4243_$1I3863_CHBONDI_2__vlIN);
 reg [1:16] _3I4243_$1I3863_CHBONDI_1__vlIN;
 cstw cstw_1393_1 (_3I4243_$1I3863_CHBONDI[1], _3I4243_$1I3863_CHBONDI_1__vlIN);
 reg [1:16] _3I4243_$1I3863_CHBONDI_0__vlIN;
 cstw cstw_1393_0 (_3I4243_$1I3863_CHBONDI[0], _3I4243_$1I3863_CHBONDI_0__vlIN);

 wire  _3I4243_$1I3863_CONFIGENABLE;
 reg [1:16] _3I4243_$1I3863_CONFIGENABLE__vlIN;
 cstw cstw_1394 (_3I4243_$1I3863_CONFIGENABLE, _3I4243_$1I3863_CONFIGENABLE__vlIN);

 wire  _3I4243_$1I3863_CONFIGIN;
 reg [1:16] _3I4243_$1I3863_CONFIGIN__vlIN;
 cstw cstw_1395 (_3I4243_$1I3863_CONFIGIN, _3I4243_$1I3863_CONFIGIN__vlIN);

 wire  _3I4243_$1I3863_ENCHANSYNC;
 reg [1:16] _3I4243_$1I3863_ENCHANSYNC__vlIN;
 cstw cstw_1396 (_3I4243_$1I3863_ENCHANSYNC, _3I4243_$1I3863_ENCHANSYNC__vlIN);

 wire  _3I4243_$1I3863_ENMCOMMAALIGN;
 reg [1:16] _3I4243_$1I3863_ENMCOMMAALIGN__vlIN;
 cstw cstw_1397 (_3I4243_$1I3863_ENMCOMMAALIGN, _3I4243_$1I3863_ENMCOMMAALIGN__vlIN);

 wire  _3I4243_$1I3863_ENPCOMMAALIGN;
 reg [1:16] _3I4243_$1I3863_ENPCOMMAALIGN__vlIN;
 cstw cstw_1398 (_3I4243_$1I3863_ENPCOMMAALIGN, _3I4243_$1I3863_ENPCOMMAALIGN__vlIN);

 wire [1:0] _3I4243_$1I3863_LOOPBACK;
 reg [1:16] _3I4243_$1I3863_LOOPBACK_1__vlIN;
 cstw cstw_1399_1 (_3I4243_$1I3863_LOOPBACK[1], _3I4243_$1I3863_LOOPBACK_1__vlIN);
 reg [1:16] _3I4243_$1I3863_LOOPBACK_0__vlIN;
 cstw cstw_1399_0 (_3I4243_$1I3863_LOOPBACK[0], _3I4243_$1I3863_LOOPBACK_0__vlIN);

 wire  _3I4243_$1I3863_POWERDOWN;
 reg [1:16] _3I4243_$1I3863_POWERDOWN__vlIN;
 cstw cstw_1400 (_3I4243_$1I3863_POWERDOWN, _3I4243_$1I3863_POWERDOWN__vlIN);

 wire  _3I4243_$1I3863_REFCLK;
 reg [1:16] _3I4243_$1I3863_REFCLK__vlIN;
 cstw cstw_1401 (_3I4243_$1I3863_REFCLK, _3I4243_$1I3863_REFCLK__vlIN);

 wire  _3I4243_$1I3863_REFCLK2;
 reg [1:16] _3I4243_$1I3863_REFCLK2__vlIN;
 cstw cstw_1402 (_3I4243_$1I3863_REFCLK2, _3I4243_$1I3863_REFCLK2__vlIN);

 wire  _3I4243_$1I3863_REFCLKSEL;
 reg [1:16] _3I4243_$1I3863_REFCLKSEL__vlIN;
 cstw cstw_1403 (_3I4243_$1I3863_REFCLKSEL, _3I4243_$1I3863_REFCLKSEL__vlIN);

 wire  _3I4243_$1I3863_RXN;
 reg [1:16] _3I4243_$1I3863_RXN__vlIN;
 cstw cstw_1404 (_3I4243_$1I3863_RXN, _3I4243_$1I3863_RXN__vlIN);

 wire  _3I4243_$1I3863_RXP;
 reg [1:16] _3I4243_$1I3863_RXP__vlIN;
 cstw cstw_1405 (_3I4243_$1I3863_RXP, _3I4243_$1I3863_RXP__vlIN);

 wire  _3I4243_$1I3863_RXPOLARITY;
 reg [1:16] _3I4243_$1I3863_RXPOLARITY__vlIN;
 cstw cstw_1406 (_3I4243_$1I3863_RXPOLARITY, _3I4243_$1I3863_RXPOLARITY__vlIN);

 wire  _3I4243_$1I3863_RXRESET;
 reg [1:16] _3I4243_$1I3863_RXRESET__vlIN;
 cstw cstw_1407 (_3I4243_$1I3863_RXRESET, _3I4243_$1I3863_RXRESET__vlIN);

 wire  _3I4243_$1I3863_RXUSRCLK;
 reg [1:16] _3I4243_$1I3863_RXUSRCLK__vlIN;
 cstw cstw_1408 (_3I4243_$1I3863_RXUSRCLK, _3I4243_$1I3863_RXUSRCLK__vlIN);

 wire  _3I4243_$1I3863_RXUSRCLK2;
 reg [1:16] _3I4243_$1I3863_RXUSRCLK2__vlIN;
 cstw cstw_1409 (_3I4243_$1I3863_RXUSRCLK2, _3I4243_$1I3863_RXUSRCLK2__vlIN);

 wire [3:0] _3I4243_$1I3863_TXBYPASS8B10B;
 reg [1:16] _3I4243_$1I3863_TXBYPASS8B10B_3__vlIN;
 cstw cstw_1410_3 (_3I4243_$1I3863_TXBYPASS8B10B[3], _3I4243_$1I3863_TXBYPASS8B10B_3__vlIN);
 reg [1:16] _3I4243_$1I3863_TXBYPASS8B10B_2__vlIN;
 cstw cstw_1410_2 (_3I4243_$1I3863_TXBYPASS8B10B[2], _3I4243_$1I3863_TXBYPASS8B10B_2__vlIN);
 reg [1:16] _3I4243_$1I3863_TXBYPASS8B10B_1__vlIN;
 cstw cstw_1410_1 (_3I4243_$1I3863_TXBYPASS8B10B[1], _3I4243_$1I3863_TXBYPASS8B10B_1__vlIN);
 reg [1:16] _3I4243_$1I3863_TXBYPASS8B10B_0__vlIN;
 cstw cstw_1410_0 (_3I4243_$1I3863_TXBYPASS8B10B[0], _3I4243_$1I3863_TXBYPASS8B10B_0__vlIN);

 wire [3:0] _3I4243_$1I3863_TXCHARDISPMODE;
 reg [1:16] _3I4243_$1I3863_TXCHARDISPMODE_3__vlIN;
 cstw cstw_1411_3 (_3I4243_$1I3863_TXCHARDISPMODE[3], _3I4243_$1I3863_TXCHARDISPMODE_3__vlIN);
 reg [1:16] _3I4243_$1I3863_TXCHARDISPMODE_2__vlIN;
 cstw cstw_1411_2 (_3I4243_$1I3863_TXCHARDISPMODE[2], _3I4243_$1I3863_TXCHARDISPMODE_2__vlIN);
 reg [1:16] _3I4243_$1I3863_TXCHARDISPMODE_1__vlIN;
 cstw cstw_1411_1 (_3I4243_$1I3863_TXCHARDISPMODE[1], _3I4243_$1I3863_TXCHARDISPMODE_1__vlIN);
 reg [1:16] _3I4243_$1I3863_TXCHARDISPMODE_0__vlIN;
 cstw cstw_1411_0 (_3I4243_$1I3863_TXCHARDISPMODE[0], _3I4243_$1I3863_TXCHARDISPMODE_0__vlIN);

 wire [3:0] _3I4243_$1I3863_TXCHARDISPVAL;
 reg [1:16] _3I4243_$1I3863_TXCHARDISPVAL_3__vlIN;
 cstw cstw_1412_3 (_3I4243_$1I3863_TXCHARDISPVAL[3], _3I4243_$1I3863_TXCHARDISPVAL_3__vlIN);
 reg [1:16] _3I4243_$1I3863_TXCHARDISPVAL_2__vlIN;
 cstw cstw_1412_2 (_3I4243_$1I3863_TXCHARDISPVAL[2], _3I4243_$1I3863_TXCHARDISPVAL_2__vlIN);
 reg [1:16] _3I4243_$1I3863_TXCHARDISPVAL_1__vlIN;
 cstw cstw_1412_1 (_3I4243_$1I3863_TXCHARDISPVAL[1], _3I4243_$1I3863_TXCHARDISPVAL_1__vlIN);
 reg [1:16] _3I4243_$1I3863_TXCHARDISPVAL_0__vlIN;
 cstw cstw_1412_0 (_3I4243_$1I3863_TXCHARDISPVAL[0], _3I4243_$1I3863_TXCHARDISPVAL_0__vlIN);

 wire [3:0] _3I4243_$1I3863_TXCHARISK;
 reg [1:16] _3I4243_$1I3863_TXCHARISK_3__vlIN;
 cstw cstw_1413_3 (_3I4243_$1I3863_TXCHARISK[3], _3I4243_$1I3863_TXCHARISK_3__vlIN);
 reg [1:16] _3I4243_$1I3863_TXCHARISK_2__vlIN;
 cstw cstw_1413_2 (_3I4243_$1I3863_TXCHARISK[2], _3I4243_$1I3863_TXCHARISK_2__vlIN);
 reg [1:16] _3I4243_$1I3863_TXCHARISK_1__vlIN;
 cstw cstw_1413_1 (_3I4243_$1I3863_TXCHARISK[1], _3I4243_$1I3863_TXCHARISK_1__vlIN);
 reg [1:16] _3I4243_$1I3863_TXCHARISK_0__vlIN;
 cstw cstw_1413_0 (_3I4243_$1I3863_TXCHARISK[0], _3I4243_$1I3863_TXCHARISK_0__vlIN);

 wire [31:0] _3I4243_$1I3863_TXDATA;
 reg [1:16] _3I4243_$1I3863_TXDATA_31__vlIN;
 cstw cstw_1414_31 (_3I4243_$1I3863_TXDATA[31], _3I4243_$1I3863_TXDATA_31__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_30__vlIN;
 cstw cstw_1414_30 (_3I4243_$1I3863_TXDATA[30], _3I4243_$1I3863_TXDATA_30__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_29__vlIN;
 cstw cstw_1414_29 (_3I4243_$1I3863_TXDATA[29], _3I4243_$1I3863_TXDATA_29__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_28__vlIN;
 cstw cstw_1414_28 (_3I4243_$1I3863_TXDATA[28], _3I4243_$1I3863_TXDATA_28__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_27__vlIN;
 cstw cstw_1414_27 (_3I4243_$1I3863_TXDATA[27], _3I4243_$1I3863_TXDATA_27__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_26__vlIN;
 cstw cstw_1414_26 (_3I4243_$1I3863_TXDATA[26], _3I4243_$1I3863_TXDATA_26__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_25__vlIN;
 cstw cstw_1414_25 (_3I4243_$1I3863_TXDATA[25], _3I4243_$1I3863_TXDATA_25__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_24__vlIN;
 cstw cstw_1414_24 (_3I4243_$1I3863_TXDATA[24], _3I4243_$1I3863_TXDATA_24__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_23__vlIN;
 cstw cstw_1414_23 (_3I4243_$1I3863_TXDATA[23], _3I4243_$1I3863_TXDATA_23__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_22__vlIN;
 cstw cstw_1414_22 (_3I4243_$1I3863_TXDATA[22], _3I4243_$1I3863_TXDATA_22__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_21__vlIN;
 cstw cstw_1414_21 (_3I4243_$1I3863_TXDATA[21], _3I4243_$1I3863_TXDATA_21__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_20__vlIN;
 cstw cstw_1414_20 (_3I4243_$1I3863_TXDATA[20], _3I4243_$1I3863_TXDATA_20__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_19__vlIN;
 cstw cstw_1414_19 (_3I4243_$1I3863_TXDATA[19], _3I4243_$1I3863_TXDATA_19__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_18__vlIN;
 cstw cstw_1414_18 (_3I4243_$1I3863_TXDATA[18], _3I4243_$1I3863_TXDATA_18__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_17__vlIN;
 cstw cstw_1414_17 (_3I4243_$1I3863_TXDATA[17], _3I4243_$1I3863_TXDATA_17__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_16__vlIN;
 cstw cstw_1414_16 (_3I4243_$1I3863_TXDATA[16], _3I4243_$1I3863_TXDATA_16__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_15__vlIN;
 cstw cstw_1414_15 (_3I4243_$1I3863_TXDATA[15], _3I4243_$1I3863_TXDATA_15__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_14__vlIN;
 cstw cstw_1414_14 (_3I4243_$1I3863_TXDATA[14], _3I4243_$1I3863_TXDATA_14__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_13__vlIN;
 cstw cstw_1414_13 (_3I4243_$1I3863_TXDATA[13], _3I4243_$1I3863_TXDATA_13__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_12__vlIN;
 cstw cstw_1414_12 (_3I4243_$1I3863_TXDATA[12], _3I4243_$1I3863_TXDATA_12__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_11__vlIN;
 cstw cstw_1414_11 (_3I4243_$1I3863_TXDATA[11], _3I4243_$1I3863_TXDATA_11__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_10__vlIN;
 cstw cstw_1414_10 (_3I4243_$1I3863_TXDATA[10], _3I4243_$1I3863_TXDATA_10__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_9__vlIN;
 cstw cstw_1414_9 (_3I4243_$1I3863_TXDATA[9], _3I4243_$1I3863_TXDATA_9__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_8__vlIN;
 cstw cstw_1414_8 (_3I4243_$1I3863_TXDATA[8], _3I4243_$1I3863_TXDATA_8__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_7__vlIN;
 cstw cstw_1414_7 (_3I4243_$1I3863_TXDATA[7], _3I4243_$1I3863_TXDATA_7__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_6__vlIN;
 cstw cstw_1414_6 (_3I4243_$1I3863_TXDATA[6], _3I4243_$1I3863_TXDATA_6__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_5__vlIN;
 cstw cstw_1414_5 (_3I4243_$1I3863_TXDATA[5], _3I4243_$1I3863_TXDATA_5__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_4__vlIN;
 cstw cstw_1414_4 (_3I4243_$1I3863_TXDATA[4], _3I4243_$1I3863_TXDATA_4__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_3__vlIN;
 cstw cstw_1414_3 (_3I4243_$1I3863_TXDATA[3], _3I4243_$1I3863_TXDATA_3__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_2__vlIN;
 cstw cstw_1414_2 (_3I4243_$1I3863_TXDATA[2], _3I4243_$1I3863_TXDATA_2__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_1__vlIN;
 cstw cstw_1414_1 (_3I4243_$1I3863_TXDATA[1], _3I4243_$1I3863_TXDATA_1__vlIN);
 reg [1:16] _3I4243_$1I3863_TXDATA_0__vlIN;
 cstw cstw_1414_0 (_3I4243_$1I3863_TXDATA[0], _3I4243_$1I3863_TXDATA_0__vlIN);

 wire  _3I4243_$1I3863_TXFORCECRCERR;
 reg [1:16] _3I4243_$1I3863_TXFORCECRCERR__vlIN;
 cstw cstw_1415 (_3I4243_$1I3863_TXFORCECRCERR, _3I4243_$1I3863_TXFORCECRCERR__vlIN);

 wire  _3I4243_$1I3863_TXINHIBIT;
 reg [1:16] _3I4243_$1I3863_TXINHIBIT__vlIN;
 cstw cstw_1416 (_3I4243_$1I3863_TXINHIBIT, _3I4243_$1I3863_TXINHIBIT__vlIN);

 wire  _3I4243_$1I3863_TXPOLARITY;
 reg [1:16] _3I4243_$1I3863_TXPOLARITY__vlIN;
 cstw cstw_1417 (_3I4243_$1I3863_TXPOLARITY, _3I4243_$1I3863_TXPOLARITY__vlIN);

 wire  _3I4243_$1I3863_TXRESET;
 reg [1:16] _3I4243_$1I3863_TXRESET__vlIN;
 cstw cstw_1418 (_3I4243_$1I3863_TXRESET, _3I4243_$1I3863_TXRESET__vlIN);

 wire  _3I4243_$1I3863_TXUSRCLK;
 reg [1:16] _3I4243_$1I3863_TXUSRCLK__vlIN;
 cstw cstw_1419 (_3I4243_$1I3863_TXUSRCLK, _3I4243_$1I3863_TXUSRCLK__vlIN);

 wire  _3I4243_$1I3863_TXUSRCLK2;
 reg [1:16] _3I4243_$1I3863_TXUSRCLK2__vlIN;
 cstw cstw_1420 (_3I4243_$1I3863_TXUSRCLK2, _3I4243_$1I3863_TXUSRCLK2__vlIN);

 GT_CUSTOM _3I4243_$1I3863 ( _3I4243_$1I3863_CHBONDDONE , _3I4243_$1I3863_CHBONDO , _3I4243_$1I3863_CONFIGOUT , _3I4243_$1I3863_RXBUFSTATUS , _3I4243_$1I3863_RXCHARISCOMMA , _3I4243_$1I3863_RXCHARISK , _3I4243_$1I3863_RXCHECKINGCRC , _3I4243_$1I3863_RXCLKCORCNT , _3I4243_$1I3863_RXCOMMADET , _3I4243_$1I3863_RXCRCERR , _3I4243_$1I3863_RXDATA , _3I4243_$1I3863_RXDISPERR , _3I4243_$1I3863_RXLOSSOFSYNC , _3I4243_$1I3863_RXNOTINTABLE , _3I4243_$1I3863_RXREALIGN , _3I4243_$1I3863_RXRECCLK , _3I4243_$1I3863_RXRUNDISP , _3I4243_$1I3863_TXBUFERR , _3I4243_$1I3863_TXKERR , _3I4243_$1I3863_TXN , _3I4243_$1I3863_TXP , _3I4243_$1I3863_TXRUNDISP , _3I4243_$1I3863_BREFCLK , _3I4243_$1I3863_BREFCLK2 , _3I4243_$1I3863_CHBONDI , _3I4243_$1I3863_CONFIGENABLE , _3I4243_$1I3863_CONFIGIN , _3I4243_$1I3863_ENCHANSYNC , _3I4243_$1I3863_ENMCOMMAALIGN , _3I4243_$1I3863_ENPCOMMAALIGN , _3I4243_$1I3863_LOOPBACK , _3I4243_$1I3863_POWERDOWN , _3I4243_$1I3863_REFCLK , _3I4243_$1I3863_REFCLK2 , _3I4243_$1I3863_REFCLKSEL , _3I4243_$1I3863_RXN , _3I4243_$1I3863_RXP , _3I4243_$1I3863_RXPOLARITY , _3I4243_$1I3863_RXRESET , _3I4243_$1I3863_RXUSRCLK , _3I4243_$1I3863_RXUSRCLK2 , _3I4243_$1I3863_TXBYPASS8B10B , _3I4243_$1I3863_TXCHARDISPMODE , _3I4243_$1I3863_TXCHARDISPVAL , _3I4243_$1I3863_TXCHARISK , _3I4243_$1I3863_TXDATA , _3I4243_$1I3863_TXFORCECRCERR , _3I4243_$1I3863_TXINHIBIT , _3I4243_$1I3863_TXPOLARITY , _3I4243_$1I3863_TXRESET , _3I4243_$1I3863_TXUSRCLK , _3I4243_$1I3863_TXUSRCLK2  );

// ----------------------------------- //

 wire [4:0] _3I4142_$1I4152_din;
 reg [1:16] _3I4142_$1I4152_din_4__vlIN;
 cstw cstw_1421_4 (_3I4142_$1I4152_din[4], _3I4142_$1I4152_din_4__vlIN);
 reg [1:16] _3I4142_$1I4152_din_3__vlIN;
 cstw cstw_1421_3 (_3I4142_$1I4152_din[3], _3I4142_$1I4152_din_3__vlIN);
 reg [1:16] _3I4142_$1I4152_din_2__vlIN;
 cstw cstw_1421_2 (_3I4142_$1I4152_din[2], _3I4142_$1I4152_din_2__vlIN);
 reg [1:16] _3I4142_$1I4152_din_1__vlIN;
 cstw cstw_1421_1 (_3I4142_$1I4152_din[1], _3I4142_$1I4152_din_1__vlIN);
 reg [1:16] _3I4142_$1I4152_din_0__vlIN;
 cstw cstw_1421_0 (_3I4142_$1I4152_din[0], _3I4142_$1I4152_din_0__vlIN);

 wire  _3I4142_$1I4152_wr_en;
 reg [1:16] _3I4142_$1I4152_wr_en__vlIN;
 cstw cstw_1422 (_3I4142_$1I4152_wr_en, _3I4142_$1I4152_wr_en__vlIN);

 wire  _3I4142_$1I4152_wr_clk;
 reg [1:16] _3I4142_$1I4152_wr_clk__vlIN;
 cstw cstw_1423 (_3I4142_$1I4152_wr_clk, _3I4142_$1I4152_wr_clk__vlIN);

 wire  _3I4142_$1I4152_rd_en;
 reg [1:16] _3I4142_$1I4152_rd_en__vlIN;
 cstw cstw_1424 (_3I4142_$1I4152_rd_en, _3I4142_$1I4152_rd_en__vlIN);

 wire  _3I4142_$1I4152_rd_clk;
 reg [1:16] _3I4142_$1I4152_rd_clk__vlIN;
 cstw cstw_1425 (_3I4142_$1I4152_rd_clk, _3I4142_$1I4152_rd_clk__vlIN);

 wire  _3I4142_$1I4152_ainit;
 reg [1:16] _3I4142_$1I4152_ainit__vlIN;
 cstw cstw_1426 (_3I4142_$1I4152_ainit, _3I4142_$1I4152_ainit__vlIN);

 wire [4:0] _3I4142_$1I4152_dout;

 wire  _3I4142_$1I4152_full;

 wire  _3I4142_$1I4152_empty;

 af_clb_5x31rpm _3I4142_$1I4152 ( _3I4142_$1I4152_din , _3I4142_$1I4152_wr_en , _3I4142_$1I4152_wr_clk , _3I4142_$1I4152_rd_en , _3I4142_$1I4152_rd_clk , _3I4142_$1I4152_ainit , _3I4142_$1I4152_dout , _3I4142_$1I4152_full , _3I4142_$1I4152_empty  );

// ----------------------------------- //

 wire  _3I4142_$1I3863_CHBONDDONE;

 wire [3:0] _3I4142_$1I3863_CHBONDO;

 wire  _3I4142_$1I3863_CONFIGOUT;

 wire [1:0] _3I4142_$1I3863_RXBUFSTATUS;

 wire [3:0] _3I4142_$1I3863_RXCHARISCOMMA;

 wire [3:0] _3I4142_$1I3863_RXCHARISK;

 wire  _3I4142_$1I3863_RXCHECKINGCRC;

 wire [2:0] _3I4142_$1I3863_RXCLKCORCNT;

 wire  _3I4142_$1I3863_RXCOMMADET;

 wire  _3I4142_$1I3863_RXCRCERR;

 wire [31:0] _3I4142_$1I3863_RXDATA;

 wire [3:0] _3I4142_$1I3863_RXDISPERR;

 wire [1:0] _3I4142_$1I3863_RXLOSSOFSYNC;

 wire [3:0] _3I4142_$1I3863_RXNOTINTABLE;

 wire  _3I4142_$1I3863_RXREALIGN;

 wire  _3I4142_$1I3863_RXRECCLK;

 wire [3:0] _3I4142_$1I3863_RXRUNDISP;

 wire  _3I4142_$1I3863_TXBUFERR;

 wire [3:0] _3I4142_$1I3863_TXKERR;

 wire  _3I4142_$1I3863_TXN;

 wire  _3I4142_$1I3863_TXP;

 wire [3:0] _3I4142_$1I3863_TXRUNDISP;

 wire  _3I4142_$1I3863_BREFCLK;
 reg [1:16] _3I4142_$1I3863_BREFCLK__vlIN;
 cstw cstw_1427 (_3I4142_$1I3863_BREFCLK, _3I4142_$1I3863_BREFCLK__vlIN);

 wire  _3I4142_$1I3863_BREFCLK2;
 reg [1:16] _3I4142_$1I3863_BREFCLK2__vlIN;
 cstw cstw_1428 (_3I4142_$1I3863_BREFCLK2, _3I4142_$1I3863_BREFCLK2__vlIN);

 wire [3:0] _3I4142_$1I3863_CHBONDI;
 reg [1:16] _3I4142_$1I3863_CHBONDI_3__vlIN;
 cstw cstw_1429_3 (_3I4142_$1I3863_CHBONDI[3], _3I4142_$1I3863_CHBONDI_3__vlIN);
 reg [1:16] _3I4142_$1I3863_CHBONDI_2__vlIN;
 cstw cstw_1429_2 (_3I4142_$1I3863_CHBONDI[2], _3I4142_$1I3863_CHBONDI_2__vlIN);
 reg [1:16] _3I4142_$1I3863_CHBONDI_1__vlIN;
 cstw cstw_1429_1 (_3I4142_$1I3863_CHBONDI[1], _3I4142_$1I3863_CHBONDI_1__vlIN);
 reg [1:16] _3I4142_$1I3863_CHBONDI_0__vlIN;
 cstw cstw_1429_0 (_3I4142_$1I3863_CHBONDI[0], _3I4142_$1I3863_CHBONDI_0__vlIN);

 wire  _3I4142_$1I3863_CONFIGENABLE;
 reg [1:16] _3I4142_$1I3863_CONFIGENABLE__vlIN;
 cstw cstw_1430 (_3I4142_$1I3863_CONFIGENABLE, _3I4142_$1I3863_CONFIGENABLE__vlIN);

 wire  _3I4142_$1I3863_CONFIGIN;
 reg [1:16] _3I4142_$1I3863_CONFIGIN__vlIN;
 cstw cstw_1431 (_3I4142_$1I3863_CONFIGIN, _3I4142_$1I3863_CONFIGIN__vlIN);

 wire  _3I4142_$1I3863_ENCHANSYNC;
 reg [1:16] _3I4142_$1I3863_ENCHANSYNC__vlIN;
 cstw cstw_1432 (_3I4142_$1I3863_ENCHANSYNC, _3I4142_$1I3863_ENCHANSYNC__vlIN);

 wire  _3I4142_$1I3863_ENMCOMMAALIGN;
 reg [1:16] _3I4142_$1I3863_ENMCOMMAALIGN__vlIN;
 cstw cstw_1433 (_3I4142_$1I3863_ENMCOMMAALIGN, _3I4142_$1I3863_ENMCOMMAALIGN__vlIN);

 wire  _3I4142_$1I3863_ENPCOMMAALIGN;
 reg [1:16] _3I4142_$1I3863_ENPCOMMAALIGN__vlIN;
 cstw cstw_1434 (_3I4142_$1I3863_ENPCOMMAALIGN, _3I4142_$1I3863_ENPCOMMAALIGN__vlIN);

 wire [1:0] _3I4142_$1I3863_LOOPBACK;
 reg [1:16] _3I4142_$1I3863_LOOPBACK_1__vlIN;
 cstw cstw_1435_1 (_3I4142_$1I3863_LOOPBACK[1], _3I4142_$1I3863_LOOPBACK_1__vlIN);
 reg [1:16] _3I4142_$1I3863_LOOPBACK_0__vlIN;
 cstw cstw_1435_0 (_3I4142_$1I3863_LOOPBACK[0], _3I4142_$1I3863_LOOPBACK_0__vlIN);

 wire  _3I4142_$1I3863_POWERDOWN;
 reg [1:16] _3I4142_$1I3863_POWERDOWN__vlIN;
 cstw cstw_1436 (_3I4142_$1I3863_POWERDOWN, _3I4142_$1I3863_POWERDOWN__vlIN);

 wire  _3I4142_$1I3863_REFCLK;
 reg [1:16] _3I4142_$1I3863_REFCLK__vlIN;
 cstw cstw_1437 (_3I4142_$1I3863_REFCLK, _3I4142_$1I3863_REFCLK__vlIN);

 wire  _3I4142_$1I3863_REFCLK2;
 reg [1:16] _3I4142_$1I3863_REFCLK2__vlIN;
 cstw cstw_1438 (_3I4142_$1I3863_REFCLK2, _3I4142_$1I3863_REFCLK2__vlIN);

 wire  _3I4142_$1I3863_REFCLKSEL;
 reg [1:16] _3I4142_$1I3863_REFCLKSEL__vlIN;
 cstw cstw_1439 (_3I4142_$1I3863_REFCLKSEL, _3I4142_$1I3863_REFCLKSEL__vlIN);

 wire  _3I4142_$1I3863_RXN;
 reg [1:16] _3I4142_$1I3863_RXN__vlIN;
 cstw cstw_1440 (_3I4142_$1I3863_RXN, _3I4142_$1I3863_RXN__vlIN);

 wire  _3I4142_$1I3863_RXP;
 reg [1:16] _3I4142_$1I3863_RXP__vlIN;
 cstw cstw_1441 (_3I4142_$1I3863_RXP, _3I4142_$1I3863_RXP__vlIN);

 wire  _3I4142_$1I3863_RXPOLARITY;
 reg [1:16] _3I4142_$1I3863_RXPOLARITY__vlIN;
 cstw cstw_1442 (_3I4142_$1I3863_RXPOLARITY, _3I4142_$1I3863_RXPOLARITY__vlIN);

 wire  _3I4142_$1I3863_RXRESET;
 reg [1:16] _3I4142_$1I3863_RXRESET__vlIN;
 cstw cstw_1443 (_3I4142_$1I3863_RXRESET, _3I4142_$1I3863_RXRESET__vlIN);

 wire  _3I4142_$1I3863_RXUSRCLK;
 reg [1:16] _3I4142_$1I3863_RXUSRCLK__vlIN;
 cstw cstw_1444 (_3I4142_$1I3863_RXUSRCLK, _3I4142_$1I3863_RXUSRCLK__vlIN);

 wire  _3I4142_$1I3863_RXUSRCLK2;
 reg [1:16] _3I4142_$1I3863_RXUSRCLK2__vlIN;
 cstw cstw_1445 (_3I4142_$1I3863_RXUSRCLK2, _3I4142_$1I3863_RXUSRCLK2__vlIN);

 wire [3:0] _3I4142_$1I3863_TXBYPASS8B10B;
 reg [1:16] _3I4142_$1I3863_TXBYPASS8B10B_3__vlIN;
 cstw cstw_1446_3 (_3I4142_$1I3863_TXBYPASS8B10B[3], _3I4142_$1I3863_TXBYPASS8B10B_3__vlIN);
 reg [1:16] _3I4142_$1I3863_TXBYPASS8B10B_2__vlIN;
 cstw cstw_1446_2 (_3I4142_$1I3863_TXBYPASS8B10B[2], _3I4142_$1I3863_TXBYPASS8B10B_2__vlIN);
 reg [1:16] _3I4142_$1I3863_TXBYPASS8B10B_1__vlIN;
 cstw cstw_1446_1 (_3I4142_$1I3863_TXBYPASS8B10B[1], _3I4142_$1I3863_TXBYPASS8B10B_1__vlIN);
 reg [1:16] _3I4142_$1I3863_TXBYPASS8B10B_0__vlIN;
 cstw cstw_1446_0 (_3I4142_$1I3863_TXBYPASS8B10B[0], _3I4142_$1I3863_TXBYPASS8B10B_0__vlIN);

 wire [3:0] _3I4142_$1I3863_TXCHARDISPMODE;
 reg [1:16] _3I4142_$1I3863_TXCHARDISPMODE_3__vlIN;
 cstw cstw_1447_3 (_3I4142_$1I3863_TXCHARDISPMODE[3], _3I4142_$1I3863_TXCHARDISPMODE_3__vlIN);
 reg [1:16] _3I4142_$1I3863_TXCHARDISPMODE_2__vlIN;
 cstw cstw_1447_2 (_3I4142_$1I3863_TXCHARDISPMODE[2], _3I4142_$1I3863_TXCHARDISPMODE_2__vlIN);
 reg [1:16] _3I4142_$1I3863_TXCHARDISPMODE_1__vlIN;
 cstw cstw_1447_1 (_3I4142_$1I3863_TXCHARDISPMODE[1], _3I4142_$1I3863_TXCHARDISPMODE_1__vlIN);
 reg [1:16] _3I4142_$1I3863_TXCHARDISPMODE_0__vlIN;
 cstw cstw_1447_0 (_3I4142_$1I3863_TXCHARDISPMODE[0], _3I4142_$1I3863_TXCHARDISPMODE_0__vlIN);

 wire [3:0] _3I4142_$1I3863_TXCHARDISPVAL;
 reg [1:16] _3I4142_$1I3863_TXCHARDISPVAL_3__vlIN;
 cstw cstw_1448_3 (_3I4142_$1I3863_TXCHARDISPVAL[3], _3I4142_$1I3863_TXCHARDISPVAL_3__vlIN);
 reg [1:16] _3I4142_$1I3863_TXCHARDISPVAL_2__vlIN;
 cstw cstw_1448_2 (_3I4142_$1I3863_TXCHARDISPVAL[2], _3I4142_$1I3863_TXCHARDISPVAL_2__vlIN);
 reg [1:16] _3I4142_$1I3863_TXCHARDISPVAL_1__vlIN;
 cstw cstw_1448_1 (_3I4142_$1I3863_TXCHARDISPVAL[1], _3I4142_$1I3863_TXCHARDISPVAL_1__vlIN);
 reg [1:16] _3I4142_$1I3863_TXCHARDISPVAL_0__vlIN;
 cstw cstw_1448_0 (_3I4142_$1I3863_TXCHARDISPVAL[0], _3I4142_$1I3863_TXCHARDISPVAL_0__vlIN);

 wire [3:0] _3I4142_$1I3863_TXCHARISK;
 reg [1:16] _3I4142_$1I3863_TXCHARISK_3__vlIN;
 cstw cstw_1449_3 (_3I4142_$1I3863_TXCHARISK[3], _3I4142_$1I3863_TXCHARISK_3__vlIN);
 reg [1:16] _3I4142_$1I3863_TXCHARISK_2__vlIN;
 cstw cstw_1449_2 (_3I4142_$1I3863_TXCHARISK[2], _3I4142_$1I3863_TXCHARISK_2__vlIN);
 reg [1:16] _3I4142_$1I3863_TXCHARISK_1__vlIN;
 cstw cstw_1449_1 (_3I4142_$1I3863_TXCHARISK[1], _3I4142_$1I3863_TXCHARISK_1__vlIN);
 reg [1:16] _3I4142_$1I3863_TXCHARISK_0__vlIN;
 cstw cstw_1449_0 (_3I4142_$1I3863_TXCHARISK[0], _3I4142_$1I3863_TXCHARISK_0__vlIN);

 wire [31:0] _3I4142_$1I3863_TXDATA;
 reg [1:16] _3I4142_$1I3863_TXDATA_31__vlIN;
 cstw cstw_1450_31 (_3I4142_$1I3863_TXDATA[31], _3I4142_$1I3863_TXDATA_31__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_30__vlIN;
 cstw cstw_1450_30 (_3I4142_$1I3863_TXDATA[30], _3I4142_$1I3863_TXDATA_30__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_29__vlIN;
 cstw cstw_1450_29 (_3I4142_$1I3863_TXDATA[29], _3I4142_$1I3863_TXDATA_29__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_28__vlIN;
 cstw cstw_1450_28 (_3I4142_$1I3863_TXDATA[28], _3I4142_$1I3863_TXDATA_28__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_27__vlIN;
 cstw cstw_1450_27 (_3I4142_$1I3863_TXDATA[27], _3I4142_$1I3863_TXDATA_27__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_26__vlIN;
 cstw cstw_1450_26 (_3I4142_$1I3863_TXDATA[26], _3I4142_$1I3863_TXDATA_26__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_25__vlIN;
 cstw cstw_1450_25 (_3I4142_$1I3863_TXDATA[25], _3I4142_$1I3863_TXDATA_25__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_24__vlIN;
 cstw cstw_1450_24 (_3I4142_$1I3863_TXDATA[24], _3I4142_$1I3863_TXDATA_24__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_23__vlIN;
 cstw cstw_1450_23 (_3I4142_$1I3863_TXDATA[23], _3I4142_$1I3863_TXDATA_23__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_22__vlIN;
 cstw cstw_1450_22 (_3I4142_$1I3863_TXDATA[22], _3I4142_$1I3863_TXDATA_22__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_21__vlIN;
 cstw cstw_1450_21 (_3I4142_$1I3863_TXDATA[21], _3I4142_$1I3863_TXDATA_21__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_20__vlIN;
 cstw cstw_1450_20 (_3I4142_$1I3863_TXDATA[20], _3I4142_$1I3863_TXDATA_20__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_19__vlIN;
 cstw cstw_1450_19 (_3I4142_$1I3863_TXDATA[19], _3I4142_$1I3863_TXDATA_19__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_18__vlIN;
 cstw cstw_1450_18 (_3I4142_$1I3863_TXDATA[18], _3I4142_$1I3863_TXDATA_18__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_17__vlIN;
 cstw cstw_1450_17 (_3I4142_$1I3863_TXDATA[17], _3I4142_$1I3863_TXDATA_17__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_16__vlIN;
 cstw cstw_1450_16 (_3I4142_$1I3863_TXDATA[16], _3I4142_$1I3863_TXDATA_16__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_15__vlIN;
 cstw cstw_1450_15 (_3I4142_$1I3863_TXDATA[15], _3I4142_$1I3863_TXDATA_15__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_14__vlIN;
 cstw cstw_1450_14 (_3I4142_$1I3863_TXDATA[14], _3I4142_$1I3863_TXDATA_14__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_13__vlIN;
 cstw cstw_1450_13 (_3I4142_$1I3863_TXDATA[13], _3I4142_$1I3863_TXDATA_13__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_12__vlIN;
 cstw cstw_1450_12 (_3I4142_$1I3863_TXDATA[12], _3I4142_$1I3863_TXDATA_12__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_11__vlIN;
 cstw cstw_1450_11 (_3I4142_$1I3863_TXDATA[11], _3I4142_$1I3863_TXDATA_11__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_10__vlIN;
 cstw cstw_1450_10 (_3I4142_$1I3863_TXDATA[10], _3I4142_$1I3863_TXDATA_10__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_9__vlIN;
 cstw cstw_1450_9 (_3I4142_$1I3863_TXDATA[9], _3I4142_$1I3863_TXDATA_9__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_8__vlIN;
 cstw cstw_1450_8 (_3I4142_$1I3863_TXDATA[8], _3I4142_$1I3863_TXDATA_8__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_7__vlIN;
 cstw cstw_1450_7 (_3I4142_$1I3863_TXDATA[7], _3I4142_$1I3863_TXDATA_7__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_6__vlIN;
 cstw cstw_1450_6 (_3I4142_$1I3863_TXDATA[6], _3I4142_$1I3863_TXDATA_6__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_5__vlIN;
 cstw cstw_1450_5 (_3I4142_$1I3863_TXDATA[5], _3I4142_$1I3863_TXDATA_5__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_4__vlIN;
 cstw cstw_1450_4 (_3I4142_$1I3863_TXDATA[4], _3I4142_$1I3863_TXDATA_4__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_3__vlIN;
 cstw cstw_1450_3 (_3I4142_$1I3863_TXDATA[3], _3I4142_$1I3863_TXDATA_3__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_2__vlIN;
 cstw cstw_1450_2 (_3I4142_$1I3863_TXDATA[2], _3I4142_$1I3863_TXDATA_2__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_1__vlIN;
 cstw cstw_1450_1 (_3I4142_$1I3863_TXDATA[1], _3I4142_$1I3863_TXDATA_1__vlIN);
 reg [1:16] _3I4142_$1I3863_TXDATA_0__vlIN;
 cstw cstw_1450_0 (_3I4142_$1I3863_TXDATA[0], _3I4142_$1I3863_TXDATA_0__vlIN);

 wire  _3I4142_$1I3863_TXFORCECRCERR;
 reg [1:16] _3I4142_$1I3863_TXFORCECRCERR__vlIN;
 cstw cstw_1451 (_3I4142_$1I3863_TXFORCECRCERR, _3I4142_$1I3863_TXFORCECRCERR__vlIN);

 wire  _3I4142_$1I3863_TXINHIBIT;
 reg [1:16] _3I4142_$1I3863_TXINHIBIT__vlIN;
 cstw cstw_1452 (_3I4142_$1I3863_TXINHIBIT, _3I4142_$1I3863_TXINHIBIT__vlIN);

 wire  _3I4142_$1I3863_TXPOLARITY;
 reg [1:16] _3I4142_$1I3863_TXPOLARITY__vlIN;
 cstw cstw_1453 (_3I4142_$1I3863_TXPOLARITY, _3I4142_$1I3863_TXPOLARITY__vlIN);

 wire  _3I4142_$1I3863_TXRESET;
 reg [1:16] _3I4142_$1I3863_TXRESET__vlIN;
 cstw cstw_1454 (_3I4142_$1I3863_TXRESET, _3I4142_$1I3863_TXRESET__vlIN);

 wire  _3I4142_$1I3863_TXUSRCLK;
 reg [1:16] _3I4142_$1I3863_TXUSRCLK__vlIN;
 cstw cstw_1455 (_3I4142_$1I3863_TXUSRCLK, _3I4142_$1I3863_TXUSRCLK__vlIN);

 wire  _3I4142_$1I3863_TXUSRCLK2;
 reg [1:16] _3I4142_$1I3863_TXUSRCLK2__vlIN;
 cstw cstw_1456 (_3I4142_$1I3863_TXUSRCLK2, _3I4142_$1I3863_TXUSRCLK2__vlIN);

 GT_CUSTOM _3I4142_$1I3863 ( _3I4142_$1I3863_CHBONDDONE , _3I4142_$1I3863_CHBONDO , _3I4142_$1I3863_CONFIGOUT , _3I4142_$1I3863_RXBUFSTATUS , _3I4142_$1I3863_RXCHARISCOMMA , _3I4142_$1I3863_RXCHARISK , _3I4142_$1I3863_RXCHECKINGCRC , _3I4142_$1I3863_RXCLKCORCNT , _3I4142_$1I3863_RXCOMMADET , _3I4142_$1I3863_RXCRCERR , _3I4142_$1I3863_RXDATA , _3I4142_$1I3863_RXDISPERR , _3I4142_$1I3863_RXLOSSOFSYNC , _3I4142_$1I3863_RXNOTINTABLE , _3I4142_$1I3863_RXREALIGN , _3I4142_$1I3863_RXRECCLK , _3I4142_$1I3863_RXRUNDISP , _3I4142_$1I3863_TXBUFERR , _3I4142_$1I3863_TXKERR , _3I4142_$1I3863_TXN , _3I4142_$1I3863_TXP , _3I4142_$1I3863_TXRUNDISP , _3I4142_$1I3863_BREFCLK , _3I4142_$1I3863_BREFCLK2 , _3I4142_$1I3863_CHBONDI , _3I4142_$1I3863_CONFIGENABLE , _3I4142_$1I3863_CONFIGIN , _3I4142_$1I3863_ENCHANSYNC , _3I4142_$1I3863_ENMCOMMAALIGN , _3I4142_$1I3863_ENPCOMMAALIGN , _3I4142_$1I3863_LOOPBACK , _3I4142_$1I3863_POWERDOWN , _3I4142_$1I3863_REFCLK , _3I4142_$1I3863_REFCLK2 , _3I4142_$1I3863_REFCLKSEL , _3I4142_$1I3863_RXN , _3I4142_$1I3863_RXP , _3I4142_$1I3863_RXPOLARITY , _3I4142_$1I3863_RXRESET , _3I4142_$1I3863_RXUSRCLK , _3I4142_$1I3863_RXUSRCLK2 , _3I4142_$1I3863_TXBYPASS8B10B , _3I4142_$1I3863_TXCHARDISPMODE , _3I4142_$1I3863_TXCHARDISPVAL , _3I4142_$1I3863_TXCHARISK , _3I4142_$1I3863_TXDATA , _3I4142_$1I3863_TXFORCECRCERR , _3I4142_$1I3863_TXINHIBIT , _3I4142_$1I3863_TXPOLARITY , _3I4142_$1I3863_TXRESET , _3I4142_$1I3863_TXUSRCLK , _3I4142_$1I3863_TXUSRCLK2  );

// ----------------------------------- //

 wire  _2I4609_CLK0;

 wire  _2I4609_CLK180;

 wire  _2I4609_CLK270;

 wire  _2I4609_CLK2X;

 wire  _2I4609_CLK2X180;

 wire  _2I4609_CLK90;

 wire  _2I4609_CLKDV;

 wire  _2I4609_CLKFX;

 wire  _2I4609_CLKFX180;

 wire  _2I4609_LOCKED;

 wire  _2I4609_PSDONE;

 wire [7:0] _2I4609_STATUS;

 wire  _2I4609_CLKFB;
 reg [1:16] _2I4609_CLKFB__vlIN;
 cstw cstw_1457 (_2I4609_CLKFB, _2I4609_CLKFB__vlIN);

 wire  _2I4609_CLKIN;
 reg [1:16] _2I4609_CLKIN__vlIN;
 cstw cstw_1458 (_2I4609_CLKIN, _2I4609_CLKIN__vlIN);

 wire  _2I4609_DSSEN;
 reg [1:16] _2I4609_DSSEN__vlIN;
 cstw cstw_1459 (_2I4609_DSSEN, _2I4609_DSSEN__vlIN);

 wire  _2I4609_PSCLK;
 reg [1:16] _2I4609_PSCLK__vlIN;
 cstw cstw_1460 (_2I4609_PSCLK, _2I4609_PSCLK__vlIN);

 wire  _2I4609_PSEN;
 reg [1:16] _2I4609_PSEN__vlIN;
 cstw cstw_1461 (_2I4609_PSEN, _2I4609_PSEN__vlIN);

 wire  _2I4609_PSINCDEC;
 reg [1:16] _2I4609_PSINCDEC__vlIN;
 cstw cstw_1462 (_2I4609_PSINCDEC, _2I4609_PSINCDEC__vlIN);

 wire  _2I4609_RST;
 reg [1:16] _2I4609_RST__vlIN;
 cstw cstw_1463 (_2I4609_RST, _2I4609_RST__vlIN);

 DCM _2I4609 ( _2I4609_CLK0 , _2I4609_CLK180 , _2I4609_CLK270 , _2I4609_CLK2X , _2I4609_CLK2X180 , _2I4609_CLK90 , _2I4609_CLKDV , _2I4609_CLKFX , _2I4609_CLKFX180 , _2I4609_LOCKED , _2I4609_PSDONE , _2I4609_STATUS , _2I4609_CLKFB , _2I4609_CLKIN , _2I4609_DSSEN , _2I4609_PSCLK , _2I4609_PSEN , _2I4609_PSINCDEC , _2I4609_RST  );

// ----------------------------------- //

 wire  _2I4594_CLK0;

 wire  _2I4594_CLK180;

 wire  _2I4594_CLK270;

 wire  _2I4594_CLK2X;

 wire  _2I4594_CLK2X180;

 wire  _2I4594_CLK90;

 wire  _2I4594_CLKDV;

 wire  _2I4594_CLKFX;

 wire  _2I4594_CLKFX180;

 wire  _2I4594_LOCKED;

 wire  _2I4594_PSDONE;

 wire [7:0] _2I4594_STATUS;

 wire  _2I4594_CLKFB;
 reg [1:16] _2I4594_CLKFB__vlIN;
 cstw cstw_1464 (_2I4594_CLKFB, _2I4594_CLKFB__vlIN);

 wire  _2I4594_CLKIN;
 reg [1:16] _2I4594_CLKIN__vlIN;
 cstw cstw_1465 (_2I4594_CLKIN, _2I4594_CLKIN__vlIN);

 wire  _2I4594_DSSEN;
 reg [1:16] _2I4594_DSSEN__vlIN;
 cstw cstw_1466 (_2I4594_DSSEN, _2I4594_DSSEN__vlIN);

 wire  _2I4594_PSCLK;
 reg [1:16] _2I4594_PSCLK__vlIN;
 cstw cstw_1467 (_2I4594_PSCLK, _2I4594_PSCLK__vlIN);

 wire  _2I4594_PSEN;
 reg [1:16] _2I4594_PSEN__vlIN;
 cstw cstw_1468 (_2I4594_PSEN, _2I4594_PSEN__vlIN);

 wire  _2I4594_PSINCDEC;
 reg [1:16] _2I4594_PSINCDEC__vlIN;
 cstw cstw_1469 (_2I4594_PSINCDEC, _2I4594_PSINCDEC__vlIN);

 wire  _2I4594_RST;
 reg [1:16] _2I4594_RST__vlIN;
 cstw cstw_1470 (_2I4594_RST, _2I4594_RST__vlIN);

 DCM _2I4594 ( _2I4594_CLK0 , _2I4594_CLK180 , _2I4594_CLK270 , _2I4594_CLK2X , _2I4594_CLK2X180 , _2I4594_CLK90 , _2I4594_CLKDV , _2I4594_CLKFX , _2I4594_CLKFX180 , _2I4594_LOCKED , _2I4594_PSDONE , _2I4594_STATUS , _2I4594_CLKFB , _2I4594_CLKIN , _2I4594_DSSEN , _2I4594_PSCLK , _2I4594_PSEN , _2I4594_PSINCDEC , _2I4594_RST  );

// ----------------------------------- //

 wire [7:0] _1I4143_$1I4488_$1I4621_DOA;

 wire [15:0] _1I4143_$1I4488_$1I4621_DOB;

 wire [0:0] _1I4143_$1I4488_$1I4621_DOPA;

 wire [1:0] _1I4143_$1I4488_$1I4621_DOPB;

 wire [10:0] _1I4143_$1I4488_$1I4621_ADDRA;
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRA_10__vlIN;
 cstw cstw_1471_10 (_1I4143_$1I4488_$1I4621_ADDRA[10], _1I4143_$1I4488_$1I4621_ADDRA_10__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRA_9__vlIN;
 cstw cstw_1471_9 (_1I4143_$1I4488_$1I4621_ADDRA[9], _1I4143_$1I4488_$1I4621_ADDRA_9__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRA_8__vlIN;
 cstw cstw_1471_8 (_1I4143_$1I4488_$1I4621_ADDRA[8], _1I4143_$1I4488_$1I4621_ADDRA_8__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRA_7__vlIN;
 cstw cstw_1471_7 (_1I4143_$1I4488_$1I4621_ADDRA[7], _1I4143_$1I4488_$1I4621_ADDRA_7__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRA_6__vlIN;
 cstw cstw_1471_6 (_1I4143_$1I4488_$1I4621_ADDRA[6], _1I4143_$1I4488_$1I4621_ADDRA_6__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRA_5__vlIN;
 cstw cstw_1471_5 (_1I4143_$1I4488_$1I4621_ADDRA[5], _1I4143_$1I4488_$1I4621_ADDRA_5__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRA_4__vlIN;
 cstw cstw_1471_4 (_1I4143_$1I4488_$1I4621_ADDRA[4], _1I4143_$1I4488_$1I4621_ADDRA_4__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRA_3__vlIN;
 cstw cstw_1471_3 (_1I4143_$1I4488_$1I4621_ADDRA[3], _1I4143_$1I4488_$1I4621_ADDRA_3__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRA_2__vlIN;
 cstw cstw_1471_2 (_1I4143_$1I4488_$1I4621_ADDRA[2], _1I4143_$1I4488_$1I4621_ADDRA_2__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRA_1__vlIN;
 cstw cstw_1471_1 (_1I4143_$1I4488_$1I4621_ADDRA[1], _1I4143_$1I4488_$1I4621_ADDRA_1__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRA_0__vlIN;
 cstw cstw_1471_0 (_1I4143_$1I4488_$1I4621_ADDRA[0], _1I4143_$1I4488_$1I4621_ADDRA_0__vlIN);

 wire [9:0] _1I4143_$1I4488_$1I4621_ADDRB;
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRB_9__vlIN;
 cstw cstw_1472_9 (_1I4143_$1I4488_$1I4621_ADDRB[9], _1I4143_$1I4488_$1I4621_ADDRB_9__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRB_8__vlIN;
 cstw cstw_1472_8 (_1I4143_$1I4488_$1I4621_ADDRB[8], _1I4143_$1I4488_$1I4621_ADDRB_8__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRB_7__vlIN;
 cstw cstw_1472_7 (_1I4143_$1I4488_$1I4621_ADDRB[7], _1I4143_$1I4488_$1I4621_ADDRB_7__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRB_6__vlIN;
 cstw cstw_1472_6 (_1I4143_$1I4488_$1I4621_ADDRB[6], _1I4143_$1I4488_$1I4621_ADDRB_6__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRB_5__vlIN;
 cstw cstw_1472_5 (_1I4143_$1I4488_$1I4621_ADDRB[5], _1I4143_$1I4488_$1I4621_ADDRB_5__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRB_4__vlIN;
 cstw cstw_1472_4 (_1I4143_$1I4488_$1I4621_ADDRB[4], _1I4143_$1I4488_$1I4621_ADDRB_4__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRB_3__vlIN;
 cstw cstw_1472_3 (_1I4143_$1I4488_$1I4621_ADDRB[3], _1I4143_$1I4488_$1I4621_ADDRB_3__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRB_2__vlIN;
 cstw cstw_1472_2 (_1I4143_$1I4488_$1I4621_ADDRB[2], _1I4143_$1I4488_$1I4621_ADDRB_2__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRB_1__vlIN;
 cstw cstw_1472_1 (_1I4143_$1I4488_$1I4621_ADDRB[1], _1I4143_$1I4488_$1I4621_ADDRB_1__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_ADDRB_0__vlIN;
 cstw cstw_1472_0 (_1I4143_$1I4488_$1I4621_ADDRB[0], _1I4143_$1I4488_$1I4621_ADDRB_0__vlIN);

 wire  _1I4143_$1I4488_$1I4621_CLKA;
 reg [1:16] _1I4143_$1I4488_$1I4621_CLKA__vlIN;
 cstw cstw_1473 (_1I4143_$1I4488_$1I4621_CLKA, _1I4143_$1I4488_$1I4621_CLKA__vlIN);

 wire  _1I4143_$1I4488_$1I4621_CLKB;
 reg [1:16] _1I4143_$1I4488_$1I4621_CLKB__vlIN;
 cstw cstw_1474 (_1I4143_$1I4488_$1I4621_CLKB, _1I4143_$1I4488_$1I4621_CLKB__vlIN);

 wire [7:0] _1I4143_$1I4488_$1I4621_DIA;
 reg [1:16] _1I4143_$1I4488_$1I4621_DIA_7__vlIN;
 cstw cstw_1475_7 (_1I4143_$1I4488_$1I4621_DIA[7], _1I4143_$1I4488_$1I4621_DIA_7__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIA_6__vlIN;
 cstw cstw_1475_6 (_1I4143_$1I4488_$1I4621_DIA[6], _1I4143_$1I4488_$1I4621_DIA_6__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIA_5__vlIN;
 cstw cstw_1475_5 (_1I4143_$1I4488_$1I4621_DIA[5], _1I4143_$1I4488_$1I4621_DIA_5__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIA_4__vlIN;
 cstw cstw_1475_4 (_1I4143_$1I4488_$1I4621_DIA[4], _1I4143_$1I4488_$1I4621_DIA_4__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIA_3__vlIN;
 cstw cstw_1475_3 (_1I4143_$1I4488_$1I4621_DIA[3], _1I4143_$1I4488_$1I4621_DIA_3__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIA_2__vlIN;
 cstw cstw_1475_2 (_1I4143_$1I4488_$1I4621_DIA[2], _1I4143_$1I4488_$1I4621_DIA_2__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIA_1__vlIN;
 cstw cstw_1475_1 (_1I4143_$1I4488_$1I4621_DIA[1], _1I4143_$1I4488_$1I4621_DIA_1__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIA_0__vlIN;
 cstw cstw_1475_0 (_1I4143_$1I4488_$1I4621_DIA[0], _1I4143_$1I4488_$1I4621_DIA_0__vlIN);

 wire [15:0] _1I4143_$1I4488_$1I4621_DIB;
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_15__vlIN;
 cstw cstw_1476_15 (_1I4143_$1I4488_$1I4621_DIB[15], _1I4143_$1I4488_$1I4621_DIB_15__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_14__vlIN;
 cstw cstw_1476_14 (_1I4143_$1I4488_$1I4621_DIB[14], _1I4143_$1I4488_$1I4621_DIB_14__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_13__vlIN;
 cstw cstw_1476_13 (_1I4143_$1I4488_$1I4621_DIB[13], _1I4143_$1I4488_$1I4621_DIB_13__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_12__vlIN;
 cstw cstw_1476_12 (_1I4143_$1I4488_$1I4621_DIB[12], _1I4143_$1I4488_$1I4621_DIB_12__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_11__vlIN;
 cstw cstw_1476_11 (_1I4143_$1I4488_$1I4621_DIB[11], _1I4143_$1I4488_$1I4621_DIB_11__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_10__vlIN;
 cstw cstw_1476_10 (_1I4143_$1I4488_$1I4621_DIB[10], _1I4143_$1I4488_$1I4621_DIB_10__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_9__vlIN;
 cstw cstw_1476_9 (_1I4143_$1I4488_$1I4621_DIB[9], _1I4143_$1I4488_$1I4621_DIB_9__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_8__vlIN;
 cstw cstw_1476_8 (_1I4143_$1I4488_$1I4621_DIB[8], _1I4143_$1I4488_$1I4621_DIB_8__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_7__vlIN;
 cstw cstw_1476_7 (_1I4143_$1I4488_$1I4621_DIB[7], _1I4143_$1I4488_$1I4621_DIB_7__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_6__vlIN;
 cstw cstw_1476_6 (_1I4143_$1I4488_$1I4621_DIB[6], _1I4143_$1I4488_$1I4621_DIB_6__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_5__vlIN;
 cstw cstw_1476_5 (_1I4143_$1I4488_$1I4621_DIB[5], _1I4143_$1I4488_$1I4621_DIB_5__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_4__vlIN;
 cstw cstw_1476_4 (_1I4143_$1I4488_$1I4621_DIB[4], _1I4143_$1I4488_$1I4621_DIB_4__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_3__vlIN;
 cstw cstw_1476_3 (_1I4143_$1I4488_$1I4621_DIB[3], _1I4143_$1I4488_$1I4621_DIB_3__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_2__vlIN;
 cstw cstw_1476_2 (_1I4143_$1I4488_$1I4621_DIB[2], _1I4143_$1I4488_$1I4621_DIB_2__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_1__vlIN;
 cstw cstw_1476_1 (_1I4143_$1I4488_$1I4621_DIB[1], _1I4143_$1I4488_$1I4621_DIB_1__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIB_0__vlIN;
 cstw cstw_1476_0 (_1I4143_$1I4488_$1I4621_DIB[0], _1I4143_$1I4488_$1I4621_DIB_0__vlIN);

 wire [0:0] _1I4143_$1I4488_$1I4621_DIPA;
 reg [1:16] _1I4143_$1I4488_$1I4621_DIPA_0__vlIN;
 cstw cstw_1477_0 (_1I4143_$1I4488_$1I4621_DIPA[0], _1I4143_$1I4488_$1I4621_DIPA_0__vlIN);

 wire [1:0] _1I4143_$1I4488_$1I4621_DIPB;
 reg [1:16] _1I4143_$1I4488_$1I4621_DIPB_1__vlIN;
 cstw cstw_1478_1 (_1I4143_$1I4488_$1I4621_DIPB[1], _1I4143_$1I4488_$1I4621_DIPB_1__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4621_DIPB_0__vlIN;
 cstw cstw_1478_0 (_1I4143_$1I4488_$1I4621_DIPB[0], _1I4143_$1I4488_$1I4621_DIPB_0__vlIN);

 wire  _1I4143_$1I4488_$1I4621_ENA;
 reg [1:16] _1I4143_$1I4488_$1I4621_ENA__vlIN;
 cstw cstw_1479 (_1I4143_$1I4488_$1I4621_ENA, _1I4143_$1I4488_$1I4621_ENA__vlIN);

 wire  _1I4143_$1I4488_$1I4621_ENB;
 reg [1:16] _1I4143_$1I4488_$1I4621_ENB__vlIN;
 cstw cstw_1480 (_1I4143_$1I4488_$1I4621_ENB, _1I4143_$1I4488_$1I4621_ENB__vlIN);

 wire  _1I4143_$1I4488_$1I4621_SSRA;
 reg [1:16] _1I4143_$1I4488_$1I4621_SSRA__vlIN;
 cstw cstw_1481 (_1I4143_$1I4488_$1I4621_SSRA, _1I4143_$1I4488_$1I4621_SSRA__vlIN);

 wire  _1I4143_$1I4488_$1I4621_SSRB;
 reg [1:16] _1I4143_$1I4488_$1I4621_SSRB__vlIN;
 cstw cstw_1482 (_1I4143_$1I4488_$1I4621_SSRB, _1I4143_$1I4488_$1I4621_SSRB__vlIN);

 wire  _1I4143_$1I4488_$1I4621_WEA;
 reg [1:16] _1I4143_$1I4488_$1I4621_WEA__vlIN;
 cstw cstw_1483 (_1I4143_$1I4488_$1I4621_WEA, _1I4143_$1I4488_$1I4621_WEA__vlIN);

 wire  _1I4143_$1I4488_$1I4621_WEB;
 reg [1:16] _1I4143_$1I4488_$1I4621_WEB__vlIN;
 cstw cstw_1484 (_1I4143_$1I4488_$1I4621_WEB, _1I4143_$1I4488_$1I4621_WEB__vlIN);

 RAMB16_S9_S18 _1I4143_$1I4488_$1I4621 ( _1I4143_$1I4488_$1I4621_DOA , _1I4143_$1I4488_$1I4621_DOB , _1I4143_$1I4488_$1I4621_DOPA , _1I4143_$1I4488_$1I4621_DOPB , _1I4143_$1I4488_$1I4621_ADDRA , _1I4143_$1I4488_$1I4621_ADDRB , _1I4143_$1I4488_$1I4621_CLKA , _1I4143_$1I4488_$1I4621_CLKB , _1I4143_$1I4488_$1I4621_DIA , _1I4143_$1I4488_$1I4621_DIB , _1I4143_$1I4488_$1I4621_DIPA , _1I4143_$1I4488_$1I4621_DIPB , _1I4143_$1I4488_$1I4621_ENA , _1I4143_$1I4488_$1I4621_ENB , _1I4143_$1I4488_$1I4621_SSRA , _1I4143_$1I4488_$1I4621_SSRB , _1I4143_$1I4488_$1I4621_WEA , _1I4143_$1I4488_$1I4621_WEB  );

// ----------------------------------- //

 wire [7:0] _1I4143_$1I4488_$1I4620_DOA;

 wire [15:0] _1I4143_$1I4488_$1I4620_DOB;

 wire [0:0] _1I4143_$1I4488_$1I4620_DOPA;

 wire [1:0] _1I4143_$1I4488_$1I4620_DOPB;

 wire [10:0] _1I4143_$1I4488_$1I4620_ADDRA;
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRA_10__vlIN;
 cstw cstw_1485_10 (_1I4143_$1I4488_$1I4620_ADDRA[10], _1I4143_$1I4488_$1I4620_ADDRA_10__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRA_9__vlIN;
 cstw cstw_1485_9 (_1I4143_$1I4488_$1I4620_ADDRA[9], _1I4143_$1I4488_$1I4620_ADDRA_9__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRA_8__vlIN;
 cstw cstw_1485_8 (_1I4143_$1I4488_$1I4620_ADDRA[8], _1I4143_$1I4488_$1I4620_ADDRA_8__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRA_7__vlIN;
 cstw cstw_1485_7 (_1I4143_$1I4488_$1I4620_ADDRA[7], _1I4143_$1I4488_$1I4620_ADDRA_7__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRA_6__vlIN;
 cstw cstw_1485_6 (_1I4143_$1I4488_$1I4620_ADDRA[6], _1I4143_$1I4488_$1I4620_ADDRA_6__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRA_5__vlIN;
 cstw cstw_1485_5 (_1I4143_$1I4488_$1I4620_ADDRA[5], _1I4143_$1I4488_$1I4620_ADDRA_5__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRA_4__vlIN;
 cstw cstw_1485_4 (_1I4143_$1I4488_$1I4620_ADDRA[4], _1I4143_$1I4488_$1I4620_ADDRA_4__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRA_3__vlIN;
 cstw cstw_1485_3 (_1I4143_$1I4488_$1I4620_ADDRA[3], _1I4143_$1I4488_$1I4620_ADDRA_3__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRA_2__vlIN;
 cstw cstw_1485_2 (_1I4143_$1I4488_$1I4620_ADDRA[2], _1I4143_$1I4488_$1I4620_ADDRA_2__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRA_1__vlIN;
 cstw cstw_1485_1 (_1I4143_$1I4488_$1I4620_ADDRA[1], _1I4143_$1I4488_$1I4620_ADDRA_1__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRA_0__vlIN;
 cstw cstw_1485_0 (_1I4143_$1I4488_$1I4620_ADDRA[0], _1I4143_$1I4488_$1I4620_ADDRA_0__vlIN);

 wire [9:0] _1I4143_$1I4488_$1I4620_ADDRB;
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRB_9__vlIN;
 cstw cstw_1486_9 (_1I4143_$1I4488_$1I4620_ADDRB[9], _1I4143_$1I4488_$1I4620_ADDRB_9__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRB_8__vlIN;
 cstw cstw_1486_8 (_1I4143_$1I4488_$1I4620_ADDRB[8], _1I4143_$1I4488_$1I4620_ADDRB_8__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRB_7__vlIN;
 cstw cstw_1486_7 (_1I4143_$1I4488_$1I4620_ADDRB[7], _1I4143_$1I4488_$1I4620_ADDRB_7__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRB_6__vlIN;
 cstw cstw_1486_6 (_1I4143_$1I4488_$1I4620_ADDRB[6], _1I4143_$1I4488_$1I4620_ADDRB_6__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRB_5__vlIN;
 cstw cstw_1486_5 (_1I4143_$1I4488_$1I4620_ADDRB[5], _1I4143_$1I4488_$1I4620_ADDRB_5__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRB_4__vlIN;
 cstw cstw_1486_4 (_1I4143_$1I4488_$1I4620_ADDRB[4], _1I4143_$1I4488_$1I4620_ADDRB_4__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRB_3__vlIN;
 cstw cstw_1486_3 (_1I4143_$1I4488_$1I4620_ADDRB[3], _1I4143_$1I4488_$1I4620_ADDRB_3__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRB_2__vlIN;
 cstw cstw_1486_2 (_1I4143_$1I4488_$1I4620_ADDRB[2], _1I4143_$1I4488_$1I4620_ADDRB_2__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRB_1__vlIN;
 cstw cstw_1486_1 (_1I4143_$1I4488_$1I4620_ADDRB[1], _1I4143_$1I4488_$1I4620_ADDRB_1__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_ADDRB_0__vlIN;
 cstw cstw_1486_0 (_1I4143_$1I4488_$1I4620_ADDRB[0], _1I4143_$1I4488_$1I4620_ADDRB_0__vlIN);

 wire  _1I4143_$1I4488_$1I4620_CLKA;
 reg [1:16] _1I4143_$1I4488_$1I4620_CLKA__vlIN;
 cstw cstw_1487 (_1I4143_$1I4488_$1I4620_CLKA, _1I4143_$1I4488_$1I4620_CLKA__vlIN);

 wire  _1I4143_$1I4488_$1I4620_CLKB;
 reg [1:16] _1I4143_$1I4488_$1I4620_CLKB__vlIN;
 cstw cstw_1488 (_1I4143_$1I4488_$1I4620_CLKB, _1I4143_$1I4488_$1I4620_CLKB__vlIN);

 wire [7:0] _1I4143_$1I4488_$1I4620_DIA;
 reg [1:16] _1I4143_$1I4488_$1I4620_DIA_7__vlIN;
 cstw cstw_1489_7 (_1I4143_$1I4488_$1I4620_DIA[7], _1I4143_$1I4488_$1I4620_DIA_7__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIA_6__vlIN;
 cstw cstw_1489_6 (_1I4143_$1I4488_$1I4620_DIA[6], _1I4143_$1I4488_$1I4620_DIA_6__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIA_5__vlIN;
 cstw cstw_1489_5 (_1I4143_$1I4488_$1I4620_DIA[5], _1I4143_$1I4488_$1I4620_DIA_5__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIA_4__vlIN;
 cstw cstw_1489_4 (_1I4143_$1I4488_$1I4620_DIA[4], _1I4143_$1I4488_$1I4620_DIA_4__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIA_3__vlIN;
 cstw cstw_1489_3 (_1I4143_$1I4488_$1I4620_DIA[3], _1I4143_$1I4488_$1I4620_DIA_3__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIA_2__vlIN;
 cstw cstw_1489_2 (_1I4143_$1I4488_$1I4620_DIA[2], _1I4143_$1I4488_$1I4620_DIA_2__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIA_1__vlIN;
 cstw cstw_1489_1 (_1I4143_$1I4488_$1I4620_DIA[1], _1I4143_$1I4488_$1I4620_DIA_1__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIA_0__vlIN;
 cstw cstw_1489_0 (_1I4143_$1I4488_$1I4620_DIA[0], _1I4143_$1I4488_$1I4620_DIA_0__vlIN);

 wire [15:0] _1I4143_$1I4488_$1I4620_DIB;
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_15__vlIN;
 cstw cstw_1490_15 (_1I4143_$1I4488_$1I4620_DIB[15], _1I4143_$1I4488_$1I4620_DIB_15__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_14__vlIN;
 cstw cstw_1490_14 (_1I4143_$1I4488_$1I4620_DIB[14], _1I4143_$1I4488_$1I4620_DIB_14__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_13__vlIN;
 cstw cstw_1490_13 (_1I4143_$1I4488_$1I4620_DIB[13], _1I4143_$1I4488_$1I4620_DIB_13__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_12__vlIN;
 cstw cstw_1490_12 (_1I4143_$1I4488_$1I4620_DIB[12], _1I4143_$1I4488_$1I4620_DIB_12__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_11__vlIN;
 cstw cstw_1490_11 (_1I4143_$1I4488_$1I4620_DIB[11], _1I4143_$1I4488_$1I4620_DIB_11__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_10__vlIN;
 cstw cstw_1490_10 (_1I4143_$1I4488_$1I4620_DIB[10], _1I4143_$1I4488_$1I4620_DIB_10__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_9__vlIN;
 cstw cstw_1490_9 (_1I4143_$1I4488_$1I4620_DIB[9], _1I4143_$1I4488_$1I4620_DIB_9__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_8__vlIN;
 cstw cstw_1490_8 (_1I4143_$1I4488_$1I4620_DIB[8], _1I4143_$1I4488_$1I4620_DIB_8__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_7__vlIN;
 cstw cstw_1490_7 (_1I4143_$1I4488_$1I4620_DIB[7], _1I4143_$1I4488_$1I4620_DIB_7__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_6__vlIN;
 cstw cstw_1490_6 (_1I4143_$1I4488_$1I4620_DIB[6], _1I4143_$1I4488_$1I4620_DIB_6__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_5__vlIN;
 cstw cstw_1490_5 (_1I4143_$1I4488_$1I4620_DIB[5], _1I4143_$1I4488_$1I4620_DIB_5__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_4__vlIN;
 cstw cstw_1490_4 (_1I4143_$1I4488_$1I4620_DIB[4], _1I4143_$1I4488_$1I4620_DIB_4__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_3__vlIN;
 cstw cstw_1490_3 (_1I4143_$1I4488_$1I4620_DIB[3], _1I4143_$1I4488_$1I4620_DIB_3__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_2__vlIN;
 cstw cstw_1490_2 (_1I4143_$1I4488_$1I4620_DIB[2], _1I4143_$1I4488_$1I4620_DIB_2__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_1__vlIN;
 cstw cstw_1490_1 (_1I4143_$1I4488_$1I4620_DIB[1], _1I4143_$1I4488_$1I4620_DIB_1__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIB_0__vlIN;
 cstw cstw_1490_0 (_1I4143_$1I4488_$1I4620_DIB[0], _1I4143_$1I4488_$1I4620_DIB_0__vlIN);

 wire [0:0] _1I4143_$1I4488_$1I4620_DIPA;
 reg [1:16] _1I4143_$1I4488_$1I4620_DIPA_0__vlIN;
 cstw cstw_1491_0 (_1I4143_$1I4488_$1I4620_DIPA[0], _1I4143_$1I4488_$1I4620_DIPA_0__vlIN);

 wire [1:0] _1I4143_$1I4488_$1I4620_DIPB;
 reg [1:16] _1I4143_$1I4488_$1I4620_DIPB_1__vlIN;
 cstw cstw_1492_1 (_1I4143_$1I4488_$1I4620_DIPB[1], _1I4143_$1I4488_$1I4620_DIPB_1__vlIN);
 reg [1:16] _1I4143_$1I4488_$1I4620_DIPB_0__vlIN;
 cstw cstw_1492_0 (_1I4143_$1I4488_$1I4620_DIPB[0], _1I4143_$1I4488_$1I4620_DIPB_0__vlIN);

 wire  _1I4143_$1I4488_$1I4620_ENA;
 reg [1:16] _1I4143_$1I4488_$1I4620_ENA__vlIN;
 cstw cstw_1493 (_1I4143_$1I4488_$1I4620_ENA, _1I4143_$1I4488_$1I4620_ENA__vlIN);

 wire  _1I4143_$1I4488_$1I4620_ENB;
 reg [1:16] _1I4143_$1I4488_$1I4620_ENB__vlIN;
 cstw cstw_1494 (_1I4143_$1I4488_$1I4620_ENB, _1I4143_$1I4488_$1I4620_ENB__vlIN);

 wire  _1I4143_$1I4488_$1I4620_SSRA;
 reg [1:16] _1I4143_$1I4488_$1I4620_SSRA__vlIN;
 cstw cstw_1495 (_1I4143_$1I4488_$1I4620_SSRA, _1I4143_$1I4488_$1I4620_SSRA__vlIN);

 wire  _1I4143_$1I4488_$1I4620_SSRB;
 reg [1:16] _1I4143_$1I4488_$1I4620_SSRB__vlIN;
 cstw cstw_1496 (_1I4143_$1I4488_$1I4620_SSRB, _1I4143_$1I4488_$1I4620_SSRB__vlIN);

 wire  _1I4143_$1I4488_$1I4620_WEA;
 reg [1:16] _1I4143_$1I4488_$1I4620_WEA__vlIN;
 cstw cstw_1497 (_1I4143_$1I4488_$1I4620_WEA, _1I4143_$1I4488_$1I4620_WEA__vlIN);

 wire  _1I4143_$1I4488_$1I4620_WEB;
 reg [1:16] _1I4143_$1I4488_$1I4620_WEB__vlIN;
 cstw cstw_1498 (_1I4143_$1I4488_$1I4620_WEB, _1I4143_$1I4488_$1I4620_WEB__vlIN);

 RAMB16_S9_S18 _1I4143_$1I4488_$1I4620 ( _1I4143_$1I4488_$1I4620_DOA , _1I4143_$1I4488_$1I4620_DOB , _1I4143_$1I4488_$1I4620_DOPA , _1I4143_$1I4488_$1I4620_DOPB , _1I4143_$1I4488_$1I4620_ADDRA , _1I4143_$1I4488_$1I4620_ADDRB , _1I4143_$1I4488_$1I4620_CLKA , _1I4143_$1I4488_$1I4620_CLKB , _1I4143_$1I4488_$1I4620_DIA , _1I4143_$1I4488_$1I4620_DIB , _1I4143_$1I4488_$1I4620_DIPA , _1I4143_$1I4488_$1I4620_DIPB , _1I4143_$1I4488_$1I4620_ENA , _1I4143_$1I4488_$1I4620_ENB , _1I4143_$1I4488_$1I4620_SSRA , _1I4143_$1I4488_$1I4620_SSRB , _1I4143_$1I4488_$1I4620_WEA , _1I4143_$1I4488_$1I4620_WEB  );

// ----------------------------------- //

 wire [4:0] _1I4142_$1I4152_din;
 reg [1:16] _1I4142_$1I4152_din_4__vlIN;
 cstw cstw_1499_4 (_1I4142_$1I4152_din[4], _1I4142_$1I4152_din_4__vlIN);
 reg [1:16] _1I4142_$1I4152_din_3__vlIN;
 cstw cstw_1499_3 (_1I4142_$1I4152_din[3], _1I4142_$1I4152_din_3__vlIN);
 reg [1:16] _1I4142_$1I4152_din_2__vlIN;
 cstw cstw_1499_2 (_1I4142_$1I4152_din[2], _1I4142_$1I4152_din_2__vlIN);
 reg [1:16] _1I4142_$1I4152_din_1__vlIN;
 cstw cstw_1499_1 (_1I4142_$1I4152_din[1], _1I4142_$1I4152_din_1__vlIN);
 reg [1:16] _1I4142_$1I4152_din_0__vlIN;
 cstw cstw_1499_0 (_1I4142_$1I4152_din[0], _1I4142_$1I4152_din_0__vlIN);

 wire  _1I4142_$1I4152_wr_en;
 reg [1:16] _1I4142_$1I4152_wr_en__vlIN;
 cstw cstw_1500 (_1I4142_$1I4152_wr_en, _1I4142_$1I4152_wr_en__vlIN);

 wire  _1I4142_$1I4152_wr_clk;
 reg [1:16] _1I4142_$1I4152_wr_clk__vlIN;
 cstw cstw_1501 (_1I4142_$1I4152_wr_clk, _1I4142_$1I4152_wr_clk__vlIN);

 wire  _1I4142_$1I4152_rd_en;
 reg [1:16] _1I4142_$1I4152_rd_en__vlIN;
 cstw cstw_1502 (_1I4142_$1I4152_rd_en, _1I4142_$1I4152_rd_en__vlIN);

 wire  _1I4142_$1I4152_rd_clk;
 reg [1:16] _1I4142_$1I4152_rd_clk__vlIN;
 cstw cstw_1503 (_1I4142_$1I4152_rd_clk, _1I4142_$1I4152_rd_clk__vlIN);

 wire  _1I4142_$1I4152_ainit;
 reg [1:16] _1I4142_$1I4152_ainit__vlIN;
 cstw cstw_1504 (_1I4142_$1I4152_ainit, _1I4142_$1I4152_ainit__vlIN);

 wire [4:0] _1I4142_$1I4152_dout;

 wire  _1I4142_$1I4152_full;

 wire  _1I4142_$1I4152_empty;

 af_clb_5x31rpm _1I4142_$1I4152 ( _1I4142_$1I4152_din , _1I4142_$1I4152_wr_en , _1I4142_$1I4152_wr_clk , _1I4142_$1I4152_rd_en , _1I4142_$1I4152_rd_clk , _1I4142_$1I4152_ainit , _1I4142_$1I4152_dout , _1I4142_$1I4152_full , _1I4142_$1I4152_empty  );

// ----------------------------------- //

 wire  _1I4142_$1I3863_CHBONDDONE;

 wire [3:0] _1I4142_$1I3863_CHBONDO;

 wire  _1I4142_$1I3863_CONFIGOUT;

 wire [1:0] _1I4142_$1I3863_RXBUFSTATUS;

 wire [3:0] _1I4142_$1I3863_RXCHARISCOMMA;

 wire [3:0] _1I4142_$1I3863_RXCHARISK;

 wire  _1I4142_$1I3863_RXCHECKINGCRC;

 wire [2:0] _1I4142_$1I3863_RXCLKCORCNT;

 wire  _1I4142_$1I3863_RXCOMMADET;

 wire  _1I4142_$1I3863_RXCRCERR;

 wire [31:0] _1I4142_$1I3863_RXDATA;

 wire [3:0] _1I4142_$1I3863_RXDISPERR;

 wire [1:0] _1I4142_$1I3863_RXLOSSOFSYNC;

 wire [3:0] _1I4142_$1I3863_RXNOTINTABLE;

 wire  _1I4142_$1I3863_RXREALIGN;

 wire  _1I4142_$1I3863_RXRECCLK;

 wire [3:0] _1I4142_$1I3863_RXRUNDISP;

 wire  _1I4142_$1I3863_TXBUFERR;

 wire [3:0] _1I4142_$1I3863_TXKERR;

 wire  _1I4142_$1I3863_TXN;

 wire  _1I4142_$1I3863_TXP;

 wire [3:0] _1I4142_$1I3863_TXRUNDISP;

 wire  _1I4142_$1I3863_BREFCLK;
 reg [1:16] _1I4142_$1I3863_BREFCLK__vlIN;
 cstw cstw_1505 (_1I4142_$1I3863_BREFCLK, _1I4142_$1I3863_BREFCLK__vlIN);

 wire  _1I4142_$1I3863_BREFCLK2;
 reg [1:16] _1I4142_$1I3863_BREFCLK2__vlIN;
 cstw cstw_1506 (_1I4142_$1I3863_BREFCLK2, _1I4142_$1I3863_BREFCLK2__vlIN);

 wire [3:0] _1I4142_$1I3863_CHBONDI;
 reg [1:16] _1I4142_$1I3863_CHBONDI_3__vlIN;
 cstw cstw_1507_3 (_1I4142_$1I3863_CHBONDI[3], _1I4142_$1I3863_CHBONDI_3__vlIN);
 reg [1:16] _1I4142_$1I3863_CHBONDI_2__vlIN;
 cstw cstw_1507_2 (_1I4142_$1I3863_CHBONDI[2], _1I4142_$1I3863_CHBONDI_2__vlIN);
 reg [1:16] _1I4142_$1I3863_CHBONDI_1__vlIN;
 cstw cstw_1507_1 (_1I4142_$1I3863_CHBONDI[1], _1I4142_$1I3863_CHBONDI_1__vlIN);
 reg [1:16] _1I4142_$1I3863_CHBONDI_0__vlIN;
 cstw cstw_1507_0 (_1I4142_$1I3863_CHBONDI[0], _1I4142_$1I3863_CHBONDI_0__vlIN);

 wire  _1I4142_$1I3863_CONFIGENABLE;
 reg [1:16] _1I4142_$1I3863_CONFIGENABLE__vlIN;
 cstw cstw_1508 (_1I4142_$1I3863_CONFIGENABLE, _1I4142_$1I3863_CONFIGENABLE__vlIN);

 wire  _1I4142_$1I3863_CONFIGIN;
 reg [1:16] _1I4142_$1I3863_CONFIGIN__vlIN;
 cstw cstw_1509 (_1I4142_$1I3863_CONFIGIN, _1I4142_$1I3863_CONFIGIN__vlIN);

 wire  _1I4142_$1I3863_ENCHANSYNC;
 reg [1:16] _1I4142_$1I3863_ENCHANSYNC__vlIN;
 cstw cstw_1510 (_1I4142_$1I3863_ENCHANSYNC, _1I4142_$1I3863_ENCHANSYNC__vlIN);

 wire  _1I4142_$1I3863_ENMCOMMAALIGN;
 reg [1:16] _1I4142_$1I3863_ENMCOMMAALIGN__vlIN;
 cstw cstw_1511 (_1I4142_$1I3863_ENMCOMMAALIGN, _1I4142_$1I3863_ENMCOMMAALIGN__vlIN);

 wire  _1I4142_$1I3863_ENPCOMMAALIGN;
 reg [1:16] _1I4142_$1I3863_ENPCOMMAALIGN__vlIN;
 cstw cstw_1512 (_1I4142_$1I3863_ENPCOMMAALIGN, _1I4142_$1I3863_ENPCOMMAALIGN__vlIN);

 wire [1:0] _1I4142_$1I3863_LOOPBACK;
 reg [1:16] _1I4142_$1I3863_LOOPBACK_1__vlIN;
 cstw cstw_1513_1 (_1I4142_$1I3863_LOOPBACK[1], _1I4142_$1I3863_LOOPBACK_1__vlIN);
 reg [1:16] _1I4142_$1I3863_LOOPBACK_0__vlIN;
 cstw cstw_1513_0 (_1I4142_$1I3863_LOOPBACK[0], _1I4142_$1I3863_LOOPBACK_0__vlIN);

 wire  _1I4142_$1I3863_POWERDOWN;
 reg [1:16] _1I4142_$1I3863_POWERDOWN__vlIN;
 cstw cstw_1514 (_1I4142_$1I3863_POWERDOWN, _1I4142_$1I3863_POWERDOWN__vlIN);

 wire  _1I4142_$1I3863_REFCLK;
 reg [1:16] _1I4142_$1I3863_REFCLK__vlIN;
 cstw cstw_1515 (_1I4142_$1I3863_REFCLK, _1I4142_$1I3863_REFCLK__vlIN);

 wire  _1I4142_$1I3863_REFCLK2;
 reg [1:16] _1I4142_$1I3863_REFCLK2__vlIN;
 cstw cstw_1516 (_1I4142_$1I3863_REFCLK2, _1I4142_$1I3863_REFCLK2__vlIN);

 wire  _1I4142_$1I3863_REFCLKSEL;
 reg [1:16] _1I4142_$1I3863_REFCLKSEL__vlIN;
 cstw cstw_1517 (_1I4142_$1I3863_REFCLKSEL, _1I4142_$1I3863_REFCLKSEL__vlIN);

 wire  _1I4142_$1I3863_RXN;
 reg [1:16] _1I4142_$1I3863_RXN__vlIN;
 cstw cstw_1518 (_1I4142_$1I3863_RXN, _1I4142_$1I3863_RXN__vlIN);

 wire  _1I4142_$1I3863_RXP;
 reg [1:16] _1I4142_$1I3863_RXP__vlIN;
 cstw cstw_1519 (_1I4142_$1I3863_RXP, _1I4142_$1I3863_RXP__vlIN);

 wire  _1I4142_$1I3863_RXPOLARITY;
 reg [1:16] _1I4142_$1I3863_RXPOLARITY__vlIN;
 cstw cstw_1520 (_1I4142_$1I3863_RXPOLARITY, _1I4142_$1I3863_RXPOLARITY__vlIN);

 wire  _1I4142_$1I3863_RXRESET;
 reg [1:16] _1I4142_$1I3863_RXRESET__vlIN;
 cstw cstw_1521 (_1I4142_$1I3863_RXRESET, _1I4142_$1I3863_RXRESET__vlIN);

 wire  _1I4142_$1I3863_RXUSRCLK;
 reg [1:16] _1I4142_$1I3863_RXUSRCLK__vlIN;
 cstw cstw_1522 (_1I4142_$1I3863_RXUSRCLK, _1I4142_$1I3863_RXUSRCLK__vlIN);

 wire  _1I4142_$1I3863_RXUSRCLK2;
 reg [1:16] _1I4142_$1I3863_RXUSRCLK2__vlIN;
 cstw cstw_1523 (_1I4142_$1I3863_RXUSRCLK2, _1I4142_$1I3863_RXUSRCLK2__vlIN);

 wire [3:0] _1I4142_$1I3863_TXBYPASS8B10B;
 reg [1:16] _1I4142_$1I3863_TXBYPASS8B10B_3__vlIN;
 cstw cstw_1524_3 (_1I4142_$1I3863_TXBYPASS8B10B[3], _1I4142_$1I3863_TXBYPASS8B10B_3__vlIN);
 reg [1:16] _1I4142_$1I3863_TXBYPASS8B10B_2__vlIN;
 cstw cstw_1524_2 (_1I4142_$1I3863_TXBYPASS8B10B[2], _1I4142_$1I3863_TXBYPASS8B10B_2__vlIN);
 reg [1:16] _1I4142_$1I3863_TXBYPASS8B10B_1__vlIN;
 cstw cstw_1524_1 (_1I4142_$1I3863_TXBYPASS8B10B[1], _1I4142_$1I3863_TXBYPASS8B10B_1__vlIN);
 reg [1:16] _1I4142_$1I3863_TXBYPASS8B10B_0__vlIN;
 cstw cstw_1524_0 (_1I4142_$1I3863_TXBYPASS8B10B[0], _1I4142_$1I3863_TXBYPASS8B10B_0__vlIN);

 wire [3:0] _1I4142_$1I3863_TXCHARDISPMODE;
 reg [1:16] _1I4142_$1I3863_TXCHARDISPMODE_3__vlIN;
 cstw cstw_1525_3 (_1I4142_$1I3863_TXCHARDISPMODE[3], _1I4142_$1I3863_TXCHARDISPMODE_3__vlIN);
 reg [1:16] _1I4142_$1I3863_TXCHARDISPMODE_2__vlIN;
 cstw cstw_1525_2 (_1I4142_$1I3863_TXCHARDISPMODE[2], _1I4142_$1I3863_TXCHARDISPMODE_2__vlIN);
 reg [1:16] _1I4142_$1I3863_TXCHARDISPMODE_1__vlIN;
 cstw cstw_1525_1 (_1I4142_$1I3863_TXCHARDISPMODE[1], _1I4142_$1I3863_TXCHARDISPMODE_1__vlIN);
 reg [1:16] _1I4142_$1I3863_TXCHARDISPMODE_0__vlIN;
 cstw cstw_1525_0 (_1I4142_$1I3863_TXCHARDISPMODE[0], _1I4142_$1I3863_TXCHARDISPMODE_0__vlIN);

 wire [3:0] _1I4142_$1I3863_TXCHARDISPVAL;
 reg [1:16] _1I4142_$1I3863_TXCHARDISPVAL_3__vlIN;
 cstw cstw_1526_3 (_1I4142_$1I3863_TXCHARDISPVAL[3], _1I4142_$1I3863_TXCHARDISPVAL_3__vlIN);
 reg [1:16] _1I4142_$1I3863_TXCHARDISPVAL_2__vlIN;
 cstw cstw_1526_2 (_1I4142_$1I3863_TXCHARDISPVAL[2], _1I4142_$1I3863_TXCHARDISPVAL_2__vlIN);
 reg [1:16] _1I4142_$1I3863_TXCHARDISPVAL_1__vlIN;
 cstw cstw_1526_1 (_1I4142_$1I3863_TXCHARDISPVAL[1], _1I4142_$1I3863_TXCHARDISPVAL_1__vlIN);
 reg [1:16] _1I4142_$1I3863_TXCHARDISPVAL_0__vlIN;
 cstw cstw_1526_0 (_1I4142_$1I3863_TXCHARDISPVAL[0], _1I4142_$1I3863_TXCHARDISPVAL_0__vlIN);

 wire [3:0] _1I4142_$1I3863_TXCHARISK;
 reg [1:16] _1I4142_$1I3863_TXCHARISK_3__vlIN;
 cstw cstw_1527_3 (_1I4142_$1I3863_TXCHARISK[3], _1I4142_$1I3863_TXCHARISK_3__vlIN);
 reg [1:16] _1I4142_$1I3863_TXCHARISK_2__vlIN;
 cstw cstw_1527_2 (_1I4142_$1I3863_TXCHARISK[2], _1I4142_$1I3863_TXCHARISK_2__vlIN);
 reg [1:16] _1I4142_$1I3863_TXCHARISK_1__vlIN;
 cstw cstw_1527_1 (_1I4142_$1I3863_TXCHARISK[1], _1I4142_$1I3863_TXCHARISK_1__vlIN);
 reg [1:16] _1I4142_$1I3863_TXCHARISK_0__vlIN;
 cstw cstw_1527_0 (_1I4142_$1I3863_TXCHARISK[0], _1I4142_$1I3863_TXCHARISK_0__vlIN);

 wire [31:0] _1I4142_$1I3863_TXDATA;
 reg [1:16] _1I4142_$1I3863_TXDATA_31__vlIN;
 cstw cstw_1528_31 (_1I4142_$1I3863_TXDATA[31], _1I4142_$1I3863_TXDATA_31__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_30__vlIN;
 cstw cstw_1528_30 (_1I4142_$1I3863_TXDATA[30], _1I4142_$1I3863_TXDATA_30__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_29__vlIN;
 cstw cstw_1528_29 (_1I4142_$1I3863_TXDATA[29], _1I4142_$1I3863_TXDATA_29__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_28__vlIN;
 cstw cstw_1528_28 (_1I4142_$1I3863_TXDATA[28], _1I4142_$1I3863_TXDATA_28__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_27__vlIN;
 cstw cstw_1528_27 (_1I4142_$1I3863_TXDATA[27], _1I4142_$1I3863_TXDATA_27__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_26__vlIN;
 cstw cstw_1528_26 (_1I4142_$1I3863_TXDATA[26], _1I4142_$1I3863_TXDATA_26__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_25__vlIN;
 cstw cstw_1528_25 (_1I4142_$1I3863_TXDATA[25], _1I4142_$1I3863_TXDATA_25__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_24__vlIN;
 cstw cstw_1528_24 (_1I4142_$1I3863_TXDATA[24], _1I4142_$1I3863_TXDATA_24__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_23__vlIN;
 cstw cstw_1528_23 (_1I4142_$1I3863_TXDATA[23], _1I4142_$1I3863_TXDATA_23__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_22__vlIN;
 cstw cstw_1528_22 (_1I4142_$1I3863_TXDATA[22], _1I4142_$1I3863_TXDATA_22__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_21__vlIN;
 cstw cstw_1528_21 (_1I4142_$1I3863_TXDATA[21], _1I4142_$1I3863_TXDATA_21__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_20__vlIN;
 cstw cstw_1528_20 (_1I4142_$1I3863_TXDATA[20], _1I4142_$1I3863_TXDATA_20__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_19__vlIN;
 cstw cstw_1528_19 (_1I4142_$1I3863_TXDATA[19], _1I4142_$1I3863_TXDATA_19__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_18__vlIN;
 cstw cstw_1528_18 (_1I4142_$1I3863_TXDATA[18], _1I4142_$1I3863_TXDATA_18__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_17__vlIN;
 cstw cstw_1528_17 (_1I4142_$1I3863_TXDATA[17], _1I4142_$1I3863_TXDATA_17__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_16__vlIN;
 cstw cstw_1528_16 (_1I4142_$1I3863_TXDATA[16], _1I4142_$1I3863_TXDATA_16__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_15__vlIN;
 cstw cstw_1528_15 (_1I4142_$1I3863_TXDATA[15], _1I4142_$1I3863_TXDATA_15__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_14__vlIN;
 cstw cstw_1528_14 (_1I4142_$1I3863_TXDATA[14], _1I4142_$1I3863_TXDATA_14__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_13__vlIN;
 cstw cstw_1528_13 (_1I4142_$1I3863_TXDATA[13], _1I4142_$1I3863_TXDATA_13__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_12__vlIN;
 cstw cstw_1528_12 (_1I4142_$1I3863_TXDATA[12], _1I4142_$1I3863_TXDATA_12__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_11__vlIN;
 cstw cstw_1528_11 (_1I4142_$1I3863_TXDATA[11], _1I4142_$1I3863_TXDATA_11__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_10__vlIN;
 cstw cstw_1528_10 (_1I4142_$1I3863_TXDATA[10], _1I4142_$1I3863_TXDATA_10__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_9__vlIN;
 cstw cstw_1528_9 (_1I4142_$1I3863_TXDATA[9], _1I4142_$1I3863_TXDATA_9__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_8__vlIN;
 cstw cstw_1528_8 (_1I4142_$1I3863_TXDATA[8], _1I4142_$1I3863_TXDATA_8__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_7__vlIN;
 cstw cstw_1528_7 (_1I4142_$1I3863_TXDATA[7], _1I4142_$1I3863_TXDATA_7__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_6__vlIN;
 cstw cstw_1528_6 (_1I4142_$1I3863_TXDATA[6], _1I4142_$1I3863_TXDATA_6__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_5__vlIN;
 cstw cstw_1528_5 (_1I4142_$1I3863_TXDATA[5], _1I4142_$1I3863_TXDATA_5__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_4__vlIN;
 cstw cstw_1528_4 (_1I4142_$1I3863_TXDATA[4], _1I4142_$1I3863_TXDATA_4__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_3__vlIN;
 cstw cstw_1528_3 (_1I4142_$1I3863_TXDATA[3], _1I4142_$1I3863_TXDATA_3__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_2__vlIN;
 cstw cstw_1528_2 (_1I4142_$1I3863_TXDATA[2], _1I4142_$1I3863_TXDATA_2__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_1__vlIN;
 cstw cstw_1528_1 (_1I4142_$1I3863_TXDATA[1], _1I4142_$1I3863_TXDATA_1__vlIN);
 reg [1:16] _1I4142_$1I3863_TXDATA_0__vlIN;
 cstw cstw_1528_0 (_1I4142_$1I3863_TXDATA[0], _1I4142_$1I3863_TXDATA_0__vlIN);

 wire  _1I4142_$1I3863_TXFORCECRCERR;
 reg [1:16] _1I4142_$1I3863_TXFORCECRCERR__vlIN;
 cstw cstw_1529 (_1I4142_$1I3863_TXFORCECRCERR, _1I4142_$1I3863_TXFORCECRCERR__vlIN);

 wire  _1I4142_$1I3863_TXINHIBIT;
 reg [1:16] _1I4142_$1I3863_TXINHIBIT__vlIN;
 cstw cstw_1530 (_1I4142_$1I3863_TXINHIBIT, _1I4142_$1I3863_TXINHIBIT__vlIN);

 wire  _1I4142_$1I3863_TXPOLARITY;
 reg [1:16] _1I4142_$1I3863_TXPOLARITY__vlIN;
 cstw cstw_1531 (_1I4142_$1I3863_TXPOLARITY, _1I4142_$1I3863_TXPOLARITY__vlIN);

 wire  _1I4142_$1I3863_TXRESET;
 reg [1:16] _1I4142_$1I3863_TXRESET__vlIN;
 cstw cstw_1532 (_1I4142_$1I3863_TXRESET, _1I4142_$1I3863_TXRESET__vlIN);

 wire  _1I4142_$1I3863_TXUSRCLK;
 reg [1:16] _1I4142_$1I3863_TXUSRCLK__vlIN;
 cstw cstw_1533 (_1I4142_$1I3863_TXUSRCLK, _1I4142_$1I3863_TXUSRCLK__vlIN);

 wire  _1I4142_$1I3863_TXUSRCLK2;
 reg [1:16] _1I4142_$1I3863_TXUSRCLK2__vlIN;
 cstw cstw_1534 (_1I4142_$1I3863_TXUSRCLK2, _1I4142_$1I3863_TXUSRCLK2__vlIN);

 GT_CUSTOM _1I4142_$1I3863 ( _1I4142_$1I3863_CHBONDDONE , _1I4142_$1I3863_CHBONDO , _1I4142_$1I3863_CONFIGOUT , _1I4142_$1I3863_RXBUFSTATUS , _1I4142_$1I3863_RXCHARISCOMMA , _1I4142_$1I3863_RXCHARISK , _1I4142_$1I3863_RXCHECKINGCRC , _1I4142_$1I3863_RXCLKCORCNT , _1I4142_$1I3863_RXCOMMADET , _1I4142_$1I3863_RXCRCERR , _1I4142_$1I3863_RXDATA , _1I4142_$1I3863_RXDISPERR , _1I4142_$1I3863_RXLOSSOFSYNC , _1I4142_$1I3863_RXNOTINTABLE , _1I4142_$1I3863_RXREALIGN , _1I4142_$1I3863_RXRECCLK , _1I4142_$1I3863_RXRUNDISP , _1I4142_$1I3863_TXBUFERR , _1I4142_$1I3863_TXKERR , _1I4142_$1I3863_TXN , _1I4142_$1I3863_TXP , _1I4142_$1I3863_TXRUNDISP , _1I4142_$1I3863_BREFCLK , _1I4142_$1I3863_BREFCLK2 , _1I4142_$1I3863_CHBONDI , _1I4142_$1I3863_CONFIGENABLE , _1I4142_$1I3863_CONFIGIN , _1I4142_$1I3863_ENCHANSYNC , _1I4142_$1I3863_ENMCOMMAALIGN , _1I4142_$1I3863_ENPCOMMAALIGN , _1I4142_$1I3863_LOOPBACK , _1I4142_$1I3863_POWERDOWN , _1I4142_$1I3863_REFCLK , _1I4142_$1I3863_REFCLK2 , _1I4142_$1I3863_REFCLKSEL , _1I4142_$1I3863_RXN , _1I4142_$1I3863_RXP , _1I4142_$1I3863_RXPOLARITY , _1I4142_$1I3863_RXRESET , _1I4142_$1I3863_RXUSRCLK , _1I4142_$1I3863_RXUSRCLK2 , _1I4142_$1I3863_TXBYPASS8B10B , _1I4142_$1I3863_TXCHARDISPMODE , _1I4142_$1I3863_TXCHARDISPVAL , _1I4142_$1I3863_TXCHARISK , _1I4142_$1I3863_TXDATA , _1I4142_$1I3863_TXFORCECRCERR , _1I4142_$1I3863_TXINHIBIT , _1I4142_$1I3863_TXPOLARITY , _1I4142_$1I3863_TXRESET , _1I4142_$1I3863_TXUSRCLK , _1I4142_$1I3863_TXUSRCLK2  );

// ----------------------------------- //

endmodule

